

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
U7hExZJod/vUi3z5N4RSr1wa48P7uP/A8O0jgaKOZBD7WNfzo6GmQd7doggkH00XJgs7nLyNvPm0
0zWCfXninQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
k253ey4kkVql4FDzRxE0SZp0nnUl5fXV3ls/4mgbh/6ghGRjfZ71MsiTZ71s3tpy77tZHD0rpNoh
xUysBr1hFwWkTjAISVTsWyokKm82DELzMzaI0lqt04f7kevY+q4XugjttAECZCOOrrnUQb5ODPuL
TN/5/7rekkgE3das7WY=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
WoA52aV8kh0bkIXA7aISXPgNn7kpio3O4wNzPv7z4wZK/v9qsQ4Fa+1FXV0tZ0D+Si1URd5Yt8PQ
TB8Mp2LGBm7aAfzTAAqLpPZr3KRYlBsnuQptgQwkquHJi1BcDR3dhZHYw2oUKeYXBoZJ80Dg1iyE
mKNc2EAX8dBe7hH745fnWjhDqr0z4schwVFz8IHUPGI/WDdrXtDdyYzuiWdux2vjC9Gao0MkqalL
zCFAkEPTT0xtWcvaccmMU2ICHf+NVjiwhEmFT/vt1jXBw7quncqpEDMuzTHteQFztMFqsgBfXXAR
/Q4rfhaHiuQ7xUCcTEngpAsL2ypgKweMgL0LDw==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Yb4xLqu3x9ghRLjHN7QkYl0tDMsZMeJQgGEQuxDwwPb+acIMCaRAm0LVh6gbF0arOSlfOKBs+X6I
1sCY01AUXvqPtXEUt+RvllN5odbTYkY9f5RujZ5aQ9olezUe3+JLEML7oIeJ23v82E3q5lEn2hpd
Yirga3+XXZGIeEC2Q5F3LdU1PK/hOr/QQAn7r3cfSPSRAYJBv2q0KFRrpHEdaRVBAVRTnMADnWqM
+83djfdVuwjO+GhXELQ+rhNH9dkL0cqvHYfgIcRG0rYfPORpbXH4Uiizi44H6tpqRpTeCgmUfW/1
kW3FxovGX7M2+iedny4BJan5eJXy8iA1/NmnQw==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pj6m4D23BtF6RtOvVlnmIzux1ocpf3A3ahzdQxUHuwpW9nlstiQd0oSmGGaiF66UD31sHUT6dfQd
yKhb6vxivgHto8LAAEiyTiUmNTH/c41wB3zGzcZFasAPOJZMvUysBGURofn88ip4eLF52/qIKVON
l8AKPEa6atmUOWXPGRix1yyvpjUnvxZ+wFAbBvP0ZsReS6AW7b6zRE+vUOJaMz0EaWEMMRdw3vLT
W/hp9Ruis3IsgHsdn6M611ZJnxSa2tuwXuWdXURUJzFjnTsi2R7EoD0bDJINDuh7T6iiDjBFdO8L
a4ER9/C3EG6IOxU+oP2sYgSHnI7dLthCIjJ+rw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
B2bb9hbJCVaDRqGS393PhTqcBLIIS3eowUvDjLX1RVvD9vYwfdlG9rjfAUVzitJwz5TOhOabACyb
mMpxy7hxgVO56ex26Ce3uZlntRRrSfXZFQT0ENioLNV+BxEHrr7uipCant7HxRFrLFt9nR5wi4m9
ZZq5zS207DucLy0jTX0=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
eqzUQVv3z3gvc1IAF6D1gFpnG3jJXG9SSewyb0B7YFlkq+2WoV55oUnb7Smo54ZcwqBR15BnF2xS
jlkL+wI6xvjzAFZaDFixez8MkTdRnrNZscyGLFWOHz7RNKwEpAxAm7RSsBEcZUaS6x+lEu8Fai/i
gBi8OQLkjYbSnKt8sfNmpRhCWxhkRR0QylraXCBqvJVR8s/2S9YSm3zj5TqvYxlJahDh9O3V0iE2
aVTZ//VjzAQrgKQboTMB5R+3O0GmOfi7O8vgrOvK/PiOq6kVyAYEvce5/1FU9VRi8AQk3Hi7BRZM
1pWTxx+bC6qDX+NQvgu8HPGpHmqeqS/CQlftQw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 506800)
`protect data_block
poe+o/1Z5OMbqSgNY7ttc2GomZFZns4h53oM6IoQWFXkR/Ys+wROz1eN3xZM0FrTD1o0+NDG6j1k
iOMxFJ7mhn5tn7QKwGXBtGBN+KGf3sHd+WzO2HF+FDgyUF7luNE0BuLc1Cc+wWKvyxICIl10w94p
DRqupypEiYrE9ehy1sg1doVWLTnlBY29HoBSaihjtRjyo494T92Q3fl+YFHF2Ar/lm5/xV9lmXdP
2X380vu91ymQD5EC5yu7LSBQiAWw9gLHkowR//e7Ce3EZMMijmB+lxl2g/ZhZ4yJ7EVWtoA9HnSk
hTcutU+a6Msc3308JwcHdn1t+SHGhJOuRa3+sl8qerteTZpmfO2o5aCptvI33IY8+6/8KwbosAsR
fEA3MSU+SV181TwkeqzE3vy1X8VWZ/jSv9M1YztwkLPml8GtMgkNGle2dKvTd1dThZeF4Y9TuYzd
yNd5/wURWmaO3X9PNzcZ79cusU62GIV3Mt5qqhbOEsspJ73BVUoNyA/t3xxGcMwQMwWakXCtzpnB
ij1Wu5UCdcJS5VnNS8JamknMVVZwovfzlhR8++lWilHGFkztKD4R9mW4ZmjpL2BPzgGzQWLFE6CI
rLFPHYY4AKCXFh9Iick56GW/WqF+9PlsLM/RzqV2dCBkvGtgGOQagIGbj0n2cYlK0+RRUTF00XrM
ZA2eiX0ADeyJih6dqHBXD1+5MbnVd3HQjO3UsEcjJTknFDhWswh1wVT6WSMYpgEsC45d2XivkgP9
2lE9Di9ewAfze8qiuVjNJQ+GUe7SxXKVgKCM0L4eVh4EB6ZEJBm+YpPWP+rjpYyooE8sWaBNfx2N
PVrfeyVo3BKCZMnCwezmE9swhiw5As5GPVijQSqm4WsxD/eUdrkrXT31Lra6HjrknANy7Kr6/iOo
JT+fhm8R3buENmKSV7RVZmyedvw+QbIIJFJo8ekY9YE4QRwo9UZlMdZSA8YnPLlvHI6U7ydS26RX
9CvwbUeIXpj/6MvLw3ObrLb31mbsDnF6dq6/3GDXT1v265rUj60ZGYhDQaPwfZo3BLUFUaOMBRH/
iv50MKvoYSGtLzAmM8hYoGxv0RtSVAKrl6qVbEmIVeySulVa1NyFpEIRRA8iBGurVIIwjTwzDdwI
KHKFTmPu+XJ1HjW61nANHQEuAmEhkr0Jcs7JGjje0NIPNsF9OfUc5ZQXOYShZTZx4FANFkDT0Fp2
eJDzX36ySeOCnwQnUFJ0p/06bJxDc8OAtzt+xZhP5v7tU07kF7oNxxl5c6By/ZpyE8sKsXoVIlBz
OgRuZr5QDq3YYOgEceUxkL57NlNjiqF9MWfAZhjjniwLC/YaLa39wF9b9s+15VVRIcCWPy0gxX98
HRO41k9Jw7M0TyfHK27KOJQygrGK4udIkEQXvvbCfTMiVxi1uw2YuGbkCcxO2W++FeHrZb1PFIj6
CAnHGY1R2gbPbvuQ9ChXWP2wxT7z39eKFHB50FhUoW+AzI8nsgdKiQSaYhtnLabPB6ztGsrxPxIE
BoFM1R23ps1dhb586OSnVnt9v8tPPEba3IB84ZLjKwL6k+5bUR0TeC42Mko0284YvnAn3AukGjz4
DRIk1aLwGcSxI1ncp2aW2PCV7UUyueQ8fCqO/vO19WpZLzwJXnKqbwAh657RzTQY0LGPJKJdt1pO
InBI9j99v82LbVLr6o3GAga+P7Lcwp8Ns/4mgQ2x9NCudmVRyjC5nm9BLKrEwovdyfUPSFIQ7ngC
eWabSuZDZG+3XRMn+PPcRZISXrQWmwTFHlwbCEFqcNxKQfA/7ksg4j1D3hTXuJZsYRMr12oNovuq
pB9jbSslxCmyNfCLTHLtATtvL2iL7LQtostAXn0P8LUKMh1VMTmLnKdjymL1Ip9kH3KGIp9lDiln
24qnZHN4q8CZ8nGjSpBrCFe7Ifwlu/yz4NzhnaOluyAaRzG7ai8Q4YPmr2u8sBLO6te5CcPGE1PV
njbxxoW+85Lar/GuvIwJUeqcWKM1CHYz+AFzABmeDPBbpZhz2hXEAJ7442mAg3TnbZVAcjUvPNoI
8jU1G38xTPdOh0AX2i0fu70e0oK7Rjrb/NCyvFu8zyiIyuwbmri/hx+dIjdN4rPA5y6TY7ZHQeg1
uUmPGQfrtxFv4kC+c99O8jpj+hg7D4vlLEEonCUoEqpXqhz4ke8qlVFQZuvMyFs3KXWnjFUbc+rG
chj00ABR1JRodU9uNSqJV+CNx7ICxIoDaxltRiy/BButdvKofrElBvpTbHCePinJfvj+VMuccXFE
q8wfnUCs3X89T8PJwUd3MI/k5jl+xm2T0z9/a+952/ploGCnN7mWL9nsyFs/7bOKK5vS9lE1b16t
WvJ+oDeoRuwfQIVS00UyE3rXCe82BtGU2E6hR1uwzM3jOfDtT8pZDhx87/9nNgbtKGJhpFSCQEa6
AaDPZmWHSYJEcLzyDBfFYZOAY4bHuWlYq9m/X2If0Gc+JjOX9MqYTVjLvKco1RHN9nLFj3eWbhgm
UFqdWhUBEFPz3zcf8rtxxcfmlCPlr9vAG32yxeHVIuo9KE8oL7wcolpH0rsDFF5RiEFMwgg0QPih
6fBLIsaM9V1AHkDyligWYyDxJmWl1GyHNbIY/yu4O9a8jXJiTYZaKp7ZbZ/1JO/ojw4YoST2yvee
6rD2rEMtcEJ201QJMnrgDtRFYmViy9zxD1kSifXFoCFtiAP09Z+HSDBYugZ+J7NnYxdzfn14JaWN
mF4q25dV1yYJAe3W5ZnpZyj8aOWuOGsCFaOj/NCrDZNkZs5e/0VJh2lDLegj+m9Sod4I3VJJXqMA
zn9LzdnjHZM5hBBnM99IUGFQllIb5pdDbPlP1bU9C4PtZIk9fVOw8AbvToT6K3xZhu9InT9psIuE
3/TBMCfmzJe/fp7xpPX8EMkPlTSPNoUQXHXDabpwGPPkgIBU7y8rFh7pbN4kaZmvSx/1z5sFSES/
qsU7LDVq/hr0mtL6KI5lT93TD4Qz7kLQORaLkszh2wG0EKkDSSx5XQtHEgy00alfDs9NctrBI8aN
7u0rRSpJF2e0Poykhn8BB0yRSYUGIJlEsEH0Dsa8QGQSR20V/vxOCHm8ZmQxjjKqAS6zTgtzkmzZ
8KVDuCvedLDnExR/rdKclOznxdg5zAccyFVeKDiBXnlghipyKPwWg+KjnjzBynGGCsxjJ1b80w4T
T52dLXq41428JDfgFGTpjXlWgzwua3TiiETJqGUPMijy3wJv21GIK/JJO3ZnEWwhr2Tjhl88XGqb
ZLurGLCpIYcV7dWGCNS2h70AnhkNL2V1nDB3tUl3QThPLpoDiPWacUbS/j1PGdh/FwDb0q1BRfqz
CC+wmR03dxO6wTDkdQ9svea3W6lTb3uFBBdi2fPdgVsgA5k38D5bj2u0ZEeYnrRPbBDhgVnm/0Gg
Q/02PlHew0YmEPe/S1IZh2VgPFGcEaOqudx2Y12OO7JVOUuAPwrJ6CgSRNPJEgz8gbPopNsQ8Xgu
r/g0GE9ZatwA1Gcwpxzfl0VfGMr2Ve3KLVwIxhHDrhkcjLDqKzBJo0Y+On2d/ejazH+bkcAqXzow
NsLCBAx7FQLDfwgUNkVaUrkfBc0HETkT1ZT/vkO9VIGn50gyl1vv97FfHax7fJeiAjDFegUWagbL
LJbcuj+Ik2kPnorOcZb4YPOlPvvgbcKbbS8S0xWiYdj2SnWWd9uUQSJIt5E+9FvQ6dEDgpLg+u2G
iqiwR7uK71vmRX9JKRreCEpJ7by4txtq6+qb85wdHMn1YwskESClaXGmQaJ9toZALQzMILEqvy+w
874BOGJeu1nX4nvs+y1lL2uTwFdEN1lfNOuGEwokio2bJDSG++LsnGlyEZDscoBt0lDdadtkDxmQ
ip552I05vphmcsGhzwn5lDTiryJj4ALohNyfUTJejKL0hJ/fGh+Sg0zE4IA7HGsL3WZkBHJn2Q2s
13r1hHjI0kYk1rdNEncoPspBL3UJEMjAzcTsdByOVatIBD0vWDFxuuw+fGkFnZOp4mFyA6TjuVAK
bBKJEubZ+WI7kUMjLK0y9OUCyHefVbY8ipWYW0yjpOf8wiyigJDNxDoQIeLxUGhr07vnX7fEQw3f
n2Yeyq1vTVb4hlL6AwpuRe/UgsLokoP5X4l3C76BjtK2jiXdn53qLbIjYblbo9Q/d9J6S7aBz8Bk
xG4v/7+pltJN4PgUzY0mH7hCd2hBk29ZW5HVDxtqanAb8vhNSvBoZDDi9/1QHMSI/Gj78N9vtl1x
cCwO4GEx4MhAxGzUYErS3R0u11yHIX6Ghd+xVDzlGKmhqc4epjQzeVVLGnPaDAK/vtd9E2S36v2o
bRyf5RhnAdzuv2RThtIVD2lUdeXpripw0e4E/ebi051iYZ6aWxv896kCSzzALDMWjS2Q4Z7lNLQu
UBo7Ra//Dudy0wAmgoqyqFgFi6d3ZeHXdunhAbJRCQnJ3mH3S3k8UchNqgcgPPiyPPcIdMv38nd8
n4VexDf2ZApvEYhhZBCj594y83/leJQdETHOL69DBbXDu5624qK5SGAMnKGqh5JdbKWv+4cBHNNk
xDzcd2i/zlBuBfU0Qe9fSSOUz4u0b5jCuds/kdrlW47s9uie7/LACFy3i3ZKPJVfYIJjoyGaU2R0
8wuheIQkbZwkToNqTJAU//tTipwlBJpqvj3jXRHVMll8Q9IKISVy1rh5dYVdf8QMT7K64TzTgGrg
rvmB+2xjoF5/Gh7p3VlTKWLrbjPYXr5npjO4YqapsHBFhV79E6N+kW04mX/bx3j6AvpjnDFdIJ1L
/1onZWbf0snkiMjRBAztCojVR+rCzRC/XGGe6GuaJjFxirHFxfWbioqpTOajUjhGF89T8XEEML8R
lha4Cu0K1xgIEIg5dA8K6JB3gZMNzKcja7He52pGCMZC5rZoPiK8NYgjboU6c+j2ApVEo+pnllBJ
HIqKJvXaqbh+6ipdIknXNXDjHdydOJJ7KJCMc0Mkoe4FKKJXrcFuBkMZipGaCkhVsAjgr6EfKOOl
59Z6i3IJwELdSbqTlSHs9E5eo8wWRV60OIL24GIFs29ti2PaHmlrlFFPsuay7MZgclEQhcOdsc+1
FpTc7VaQdipa/+jrp3GDUC3MhrDscIQJMtcApWSZ7ZWW0NKWhki3Weo7MvfLg2RBT7dmZZqhrzdh
GJDc2sOtS7quRVCvuxAr8rG14a0/wFBGsqMLxGnRLK4SOUPKGJuRQ/kFJs97oWXvOO1smMohxdBP
R8vKJRC+T36xwUYBA58kI8q93K3yZ7IUOp7yaB6CzHY4v82iomWr0y000Na1GU9B+6Z5FmE+5/bh
CAyx7c3FfIMha1JNin4WinAqF7aY3W66uLUIWmdtjaX0xiOXODqL/WBJ0dY2vxcznoVGmS58X2IE
Fmrj5m8gdZ5y9Mpf2BAO95U2iAWCIi3vjZ81S90Pdwbf0pPt4odES646NoY1yIOdXMW5lgNSP/Un
EAVqtqzad017/wEbz8mXcq3I5BYRWLRMoC2azY0mIX0JW0xuB1OuB8ugzyV5nK7DW2dTiNfKmEl0
PlFQ/8Ve3w40wgeOYpKbVOWQOVE8PmsijF/471yFq6x/0rhhOZ6nR4A2PA8xzAA70dqfMgFM9lru
h7aS5Buvt82UIfQboIX8mSeUieo8a/61mjbAq/cvdJ6trZkpCZbAIVN8YjoX4OAT4gu0/gw27fxr
K6kvIEvKIHt+syh2hEFmuF/Gf1gLo2HA805p+zsqUN/fLGtRz8mWLnt0JXtbuISJH86cqtA1RJaz
qWsnvIldVqBrdsamrnv5x7Y0lL/QacFOuW7c2MoW9Uy5X4ANPngEsQa+K5vlD9VyCP7pRDKdATuJ
ZJnGAmKm0pXGeF4nnZ/vyqDI6iUxm1NkYUl/7tBxBBWmOJRpF5GAQPjwvEVMPOlv+c1C6wrUqWbF
Uzjv0mGXIduG91dq762B0yExDX2UEGBECdtJ2O6qNB91ZzcN9GvB0iILqpiXmyNBni5lv/Cq5TI8
M0QFG8vMS/kU4WJUdLB/JUsALAc+2WOxYRJCXF0prTX5LmAFpH13nCGpN68EXcJbOk7q5pk5+OOk
zeCEP+RJle5vGt73tdmpzdpT9eSmCPJk40CDzOBviZp9fruL3BWf1/adRz2IHUbBQby8gGn2lI2x
sUnZcngONOo9jQ2xilMJEiA8aZsGCx3AHZwtDy5AstmiImGBqSYLpd16/QNcMWpmGubSs0F4aRK2
aqL2t1ffgzYDAi1qMgWy5UIcWwwGDSEDPi86ArEFnAktKPFF/rQa+86V+MVEKbEI1+x3qAiVu9dY
GvCKIfVZuLqEWE2teLvHgmET3pXrTwywYRzb71PgBAi3zF+3KgmJBnFBgyk8mAKOY93tNcZN6x1V
dq1OhX5rJ6ncTve1vZCnL28U0ffWSYw8v+BNDf/GYq+Tus6qLFp1GCwe2VKwl5sk2VJrdo+4/Eu3
2cWLCImbOzic/WHFvI889zJD76wnztHoIr4gYSo7Xh4y6u+wRP7Nno704YpxXZYJokD0D9svtagb
EzbtNz1ZSdwRAkfGMElsC+7r0ALmBbm5YtySn+ZCNXz41vK126SN7ojKEi3axER6C8LRs2C1CvHe
3q7acRG5EdNzHWbcwpI+wCpZKjvdG7LDRQAydX2nGvh8/ZuSJTB0zuJ7JVyZi9UK2ySBkkjKbfFw
ar5DmuStdo9+ARSJTv6wjEzIYolY7/0nehPWCBAp54UsEFwM+p1ZYJOAstNSUZ85k3Gow9H0vAFg
5aWUx6zxU6z2/rcPDT2EdTWsynJ4VVvw5Qm0ueaWL9NlIjeGhYxUdf9Zyxi4b0dYyRhxRY7ODJEQ
OLz4gyRDYyJRYnkEx2vwWwe/RUqLNtA8mVeS/2ycpc8mdmcztib8BkLg5AOZDdN1rNLdmy3iX3sR
OfLmo+MgfbJSwnfYdStATWsChO9vKACkxyV/0AsjQFzirQOmxz/b92zxuk1GtOOnaR0at+3NXgnt
0n9TJ27WFr2lMQG1vPy4yEuosHqDTmCsSSblxw7zDyyMyiJYxpDjnAFSadVQQHX9v31zpJpAB1WV
/WUtjPRi1Ocx+x8oFjmk1NrANq+PK/6jMIMuMTJ4/fb9RHM3DsVWF6QxwifDFRin4Ync54RaRaZs
62k4JOhmuxynxa6xGi7YSrOvkc3Zk9s/iuDSsv5nPOzb2uUPuOBZYVnam770zhimvSS4u1lEK9rZ
FJf+MB5L6H6HHS9L+aJ4GD5XGUSGuqoGb+LzJlNEVvfOfixzZPa+QbUb5sO8JjZTv+eL6tuAkK4y
4cDkhX58WgTg+IC/dSQu6Euu4uUQXXOcRfMOeoqBJrhnzx/XsPD2ciS3Ndp3CDrDt2nqjMQgkFlr
GZ7k6n8micoru42sEEJuL3nf4fmnN7ryq7XEqGNC6JrC4cMucWjbU29JK9k6ZiH9Put5R04rxMcF
C0bYkg/LV4eTHewD5HPDyS0jG71nRmkA7pIGCf4MtJ+KYeNwoR08/VvxUHepJ9KTCyDzrgVRh/Xj
prIM9gqyxkMUt39ZXt+gkW0RGy1ZgpJDDjC8n15h3Rsbwk/Vp2dWyiQcZV36jl4/EjmAG4pkZi8Q
Dl7OWFnZc53Tw8XrKyLvTumKctQIVhNsG/Y0rQlr/wvveoR7tZ1HxE+KYPdxtfdvEm66PwqeMTKC
xzjVRQLVNX0kVHAXMOdF0zyNsRPI/InBdNOrEamqGEGqu/c9Oa9jXYB6CcMyYlnC2M5/X7SInUsB
NhU0K5YX05YcJAltwhT8waJ9zLv2xTnF8WtA8hGdotjN5OL2+97MyLdIO/XSEE8Mbn4gHRwnK1m/
isa4SpDYqhbRIaHu+ef9jd/p70IS+thyQOXMOcXd20W+j4JEwfDizAGEa+Na+O0gRmXFIxXl6c4T
1NRujiPnXfAblqu4uUhZsWdPeWDRUGGceshQvaLrAvMnjXtswIOHHPVs1tV5y1t3glUy545bDI9u
UdALzKg4kuz2vO0tZE8hxHeudpPR7Ju2blTVeBaAWCr72Xi9LierJ8Isu6wv/BWPgXyi1aELcM1n
W3OaULSdZtqaBczYGC+Yht/ptYnqf33xP4/FYGFUfyT+NnuKjChZeGMZqIMZQYO2dwnXtFMH/UEQ
yWmK6N5bu0O7XY3TBrI1Hc0oiNXx+mNJBlHYSmQOD/S/O3D/M/zYh4Al1ZlZqnmNpyTqrKsrnp/H
ipNbXp4V3wnVzfr0KObC8qB2Ks1WZnKJBcRkdlf7dvzbYfns8a/PVCbpI/hhecbhQ1xbOnT3jAfe
FUR8RcQu5OwsQSFcZuYJ/eFvk6w4a6b/wF0Ev0v5npfGzaJie+pvxMRhCnmnYG+vupTDGjnwrSX2
PvQQfynZhK3KKJ1sbHYUuw2V2Eca6i+YeIqELkWlx7AeClG12v7MI5Y089Bii2CG7JeYZ+eDe/ZE
0PBuXmH1ORaPUX3QmPXkk5qeJy9X0OMyRLF1GlTLexES9iT4vgPAKA6K/4PvU0dPzIr2wP3gYHeK
whk1gnFImFg37BQrUbRELXY/3AqNItvklxTFs/KaoW2iVRC8Et0YC8fEBK+fBBgp+d15ZZX4GBqK
ffgkzfvEEtVRphB8/iyMCxGL1RTpYwEAlXZUYG4Md0L99jTuLSwafWeaznuHvzBu2IW/HWIr15L2
HlIu4lgAenA5HfpCcxA2IEarpJFIlKHmJ0gLJPyGkXpEapXQr1Pz+Jg6FkV6tqj7kzRE78OF2wAj
iq8wC3bbVxm3ZELme4fC/4E71GCVCs4JrUmkT/ZsVdnl7aSeO2BwJvzDn7tBdQiJJXRq/5L1ZQEn
UH2voQTrYdppjH7IbFpm5adMtt1gqdsFI6s9K+eO6yE9vNuIjhGr8wewfZQtCTIIzwmvtSP29YHf
zovADfsR8tF2W0niT6DveLd1EbWJdoUs4SlcnWxLpCfYIIOyRAMPGa0I5OSXzjhYRnOiY1sDrBNl
c362x99uvdfi6658VBN+DkBxKG346xeQX5OHCfPTP50w83dTrj1zJlb6Xrs0UZM7/z9ruemGl+LF
X3b4jnAl6zf3yXOh2aMh4z2XspDZzkC4qW9IK4umxqonOVuSoF6TpC7w9xc9larRxHwGExUAto8b
Nx3IX1E8CGbURZo5jnqB34kmLiDwpWrTzCEMoXoH19x8WaoQ1yRkT/8zcWAspvokV+kbFQwHpWTa
jxh4TbIJseSyYC7dACtXSI4kdnrXXqCTCAdJGCSsf4+rr23lzqjzZvML+J/FXawHSgTEStLQviJS
qq2F5T7VUwW8J9IXcy5f/w9Roa8wPcnw5vs6f02I/vMBAYDDYkBeSLZY5LQvj47WyG6H5FHm9lM5
eRxAGMSqPKv662oxDZg65m3FXXroE4CBkdT2PTFPM35ZlC1em5TT5AW9vZgELOe37aQiynbVfnI6
kr1CqrqZBQgydw/dj3ZgaJOj7U92lDr/wQZyDBlWh1yUWNzuLktamKFWmwdyjD4FqFCJV02YnBUX
I3wU+PVlZBpfxozDHfyVImz3AurgnWcesofgVFYtrx+Y9qbqKHaECLUpEvP8egzrdkGt0bbHa5mX
0gI3yetBU0/6jIWDaJmKARmOTWt+oMgcsMbE/kD3zzw95b6xpJaV818nUJ/FJvjRkPoezkj5SGJW
Bb8hoJJL717i9nZIs86ElR/fFftpuMZvyAINWuKClbEgJ+KZAnTFyVISZiPEmc5WF7jRo6QX3Lvh
oM+qD1oHmczy8Ytkg6lw4s45gTA0JTxtZ2jlubtUizGwMhwACZxVt5OdmzDyVqIMNj8YL3S7srXm
GSUTN8F45dGGUHZ/jkM9e4qocxBkGb3EwBJqRgBz5qDY/f+x6RQJ9ctxt5cXOVY/+l1m9q42V8+j
NAFIZH7v5eP6uRsRIgIv0hpi+qdqPUX4MvcHn3nbkXjMTF9hWjXyNftrKhqtflKwE8oToBl6eG57
geq8wr7tCH/Tx//pU7vkGj0R0INkrIEbspj3uMipzAl7B4WlqDEurpYmGnK+UsY3iS384IdRMieX
eO034UX886ZsF9jZMJyWe4BZnBezsfWVzHbhgf+c/YFTy+946bYvCIpnbqmCDsscAtPJXuj3rPT4
3boJPQlK9QchCyxtiKqTJc2l+Hq4Zl8XuCnYGuGac3WRI9+HvfmKXh9zSlX5JAeHNm7Xn8IMgedb
PkoHUrUJ5MvpB8IjgxhckPuZo+zz/szC/vyVPYUJwOs2coxeHfaITGqXHswShQ7xD4JQnaj1MsKT
uxBOksyXRqszjpQWz/ZWFLnYHExNEh/DvGR0ycWHAnV3ac1PLp9Cf35WLj5XxLoOd8Iu2unJkJbp
Au8p3IHX667ISMx1XUyrZBjP/QjvsmjT2u2LJDN6QDzlJhRMoR71ex2sUaR4nea8CXuWNLVxwmpR
PdgpyfwO3o/P6ZtkTShyolrHZXcPuhZ7++9MPQ1xNRmMkYHWcuAGvqLzDk8NHEXNPEmXW6jt1IKR
KfFRWusVcFyFkspTAT5nJb5r3TnQvN/lLJ/F7AUgb2JOjnYIvGtBVO/Ttc4vsJlkbROncy/8JPqk
COuACRS0TwKXps91QnL20rOtxmuTFdPSby/dpKI9tbKt00fKYMsOWxwyqQCCsinitpGXWN2js3PF
/13z+pfVdq9sMby9xKW7DGrG810PGbQVMhS64m6QZMcbTPjEIhrggyBSgCssEp1wv4Xg7/wSWMc9
Gq4uC8P20/6G5ed5ZqPMsurfqdbqPAmImMaxkQFRCnuyAbShUZz02frYssUF0iGAYQHC3zUQRkOv
Exqo8NmKGvzj+17b7254g569NL+Xb2iiuJg+eDodRI7js886WhTZC8F3YCfM1j1NO3xzx3LROTLn
oExk/3PXK8QLe63640g3hsTk6x/P42t0f7cGk+HetDqH7ia15UUVuBGbObDqKVpE3wDdp2goAGhb
HJrnh/e2pxmAMqC3wc302dcOyxNTNWlWjdMN79JtYdOSsnQ89jn6qeeEBN+tF3NXGLblBZK4CvCB
x/GRjWc3v6fJDAmgUhz8UQUQw/9RtnUezigNAK12Y2KAosH02dCERTgUgyXKVwB7CY0LbXRw6ut8
zdFjv+gW/Ukge3+RKwJL1QNx2NpzN0irZdGmbjymRqsSah4HqkDDamkA6/ZvYkwpFa828xxnR4if
aeB5GPU6uRwVl/+bVtviLyWY3Tf1qZ8NrvWVQJbL2i46KjJiO1jLbfxXaz1Gnk7PxDvoC63Arlqm
0mShT8BW1YIme13Euu81NM9+YaBTIhFjqoEz/BtJNYmTXutipgO5MsF77S0cRkXBkP6Tq7H/JjdD
ZnuI0NYGheZOkurYkmiUr2nhda33ih6ePYv3WmT5/XwWBnbqCDLTxHxaaweGJHpgecjrflRatM7p
GEMOPmZzKb8ZVzWwk9j1hk39bcXjih+SpoWYVZKdYnJ6+n757k1QT+UTFUdkWdufxXDbrxRVJaz2
hNqHKNWsNTf1QTwcgsf5IPtpOAlc8GkSdf42n8cXX7mDYSBx2Dl0x3Gh/x2U4ZVMBdmONBEjBW59
C8cA/0DulhTCZqQKi3/A1X9Nh6vaEeB6CqjbuLhr/AUA1+gryLSp5Y+crVjjpjTxcnIe8minrq5l
tgfKhAFzXVWHUhU/PxVngxe5qNcNsUUtyj6A04ClCzZxHRAgOO8VJRqkHgocHEL1kWoIOMZ6Cq6n
qnSgwanpqD0tHoNSXQUS6HLV8UtEn7zLkAbQN0AUYcxNhLFC2sSfmAim9qaY+M4y75oza5Gt8t4q
BiJJec9CjLzz3dIuuDWgOTlfH259O5wcEqxdxeQe1RRHCeUQtnDhAAqoF5a2wmcZg8j4oQuBAyay
Vo8iwsm3ByhG78PL7ArgakB45PObp5G8Mzr0ejUiRVaXiaMWvmdzPxt++v3M7ztEoUgnjbH9vwAA
NQXH84ggJo2RElwnUmnRxnPII7bcvDu6YpZlnfyAUQ6VYokZ6LkSyysBtsKnSi/yb6YyeqrVmHcm
pY0P+dSiZKMGM145LWv1fOyetstkeklrPzV4MRRFsLkgiYTWHGrL/mUYaWH7m9NIfoIOibS263jz
B2vRDj1KsnUYCtkjOQafY8EQ6yDpZiJRVktgLrRcVJykAURNcmrKh7Nb0yZ2xu3218fd/Vlxgvea
4hJ9rSPU0NPmWCbeeWrs9YxSB0aeFKp4kcjfjh836wyvtUX+03P89n/TlMiMojboKwm7mPeJB/yp
uDDQZjJPy2sTrcT8QDCKtCO0bdoCI/RZoRN1A7iN4P0SiQYEVRUFzsH96kItc7F56vd1r7jhApG5
ZUMtUQaq6THyNtKNlCpjh3SZfUHFrx8AvRQxS+Rg6NJQ4XB2WHKuQ9iApQViw/y9S0NYX5a6/hB/
9Thvn0oXJgvQl9uMKWymJrOe6/xGfTzZ40TCzGYfKCR1+lvX7J4OnGCnL/g6as2WmTKaiQmFS0wa
QzLHwjuPYcD9nJKbsS5Q30/cO4LeiIkkRsqA1b6R+Zb0hEsLD/He3zE6JdSLQQRKQt+6e34XKuao
cMQSGudBcH8AzhS79R3DFc1OarWzRE8AqN1hyO+Cmf3pGWhgP4KSCO6HdtkpojasJliNfBPRyrLE
yA5Ovh1N9ujoN2GOhnIv84LD2HAkj2AU8Hss5Ij5lENXelwYAUYIQjFJ1KgQyMvx9Rn9IBEKCSH6
HGNcoQfKHvhxQQ41v/rGHuJN1UTnTPmz0QudfqQVftqLDMozJsWKebIkVSttYEJ/WKATE9+2Q7cc
DKzsy1RSqlhoLhY5qeV2FAGqL4UjoNkm6E0uKRhNTmhkPDFCTkvxmiNdEf0+Uhl0OFO2Ykvyb8SS
/ys99cHsHhZQzNGZvPSQBm85AzUpyVbkUxtVW1Kfns5YkUeIAJC6S99c6QmNH47kLSmgKhN6Kt76
fLA2NBzj75Iyf7/1qTRjUWdfyCzQlvCZmwCoBUyvFoPm3+YtEsmTCWenSt7ICbMQEI2PDfUCfcR6
3vgq1rjuLqQ8ZojbF1G/4lymhKmVoA5kKijSbTDen0G8gG0RgiOnD73dfY8vKjOLjK1NdRFacXLQ
i70G4Uk6LbutJ5eXhHDB31bnRYnkP23ISrhZTDDvlsHVcW8C1lmq9eOpTaM6YvATKTfwxdJr0ogj
2Lpq1ejmFvd8k/xphy7z5wIi+67Wq3ZodzJgekdIFsmeYLHX7kmS0/seIntKqRw3Y42Fg9p3Bqcf
i6W7zUDlziJ4fv++UtoDT6424LMA2klOtSIXv+011PnaOjGPvDz8pe0hIgdPPGndcsC5ZyX89AMo
xE00dQYuaPECvJWE6sJqzlkuz3z0rKSi9oBp+kMzlgd0Zjj9eleQVS0G0GLCylfQ8k9syfsl2DIq
ik82HQ5KM5h7l1dvntM9u2F434JQvQVbI2pzkas/8bfM1VqZw9ftbGNmo6uasUkRwh3B4Y/P3T1z
ZYaz7nyzL1IyQxu1AV8fHYRqg2ikfmADeIs1DDZa6PhajYrD0iM9TFUY321uXSuu72zTiYr4ElEc
RY4m8NZJ2C5rKOegvE+wg0rsCE3YEDiSMqxbkr+2v417EAF5JvcPv/EyTrRnwgunzb3/oqDsjzc5
A2U9oithpIzoAXxiQfI3G+uWrr1LEljCtOjng/UoRx2xqFhvVFWcHHEfAcGWcz2lAittVUpDhQ4j
+Hwb67bY/aYH2htrbiGALAXSzZ9IRh5gYQmL+gw1C7UydzQjXfYZK+15JO7nsQqkyVAA0Cdk2WL/
wMkh8TgUQdy4dnJhuodufrEsVWPm72eM62PKQsFRJERATUTcN8305EslEAA/EaNtNYflA4L2bWA6
oSDMG8DDwTVuUyuVoKNp7m+qDi9EFoTfs2aCXMQFADUQXlk/nVQvfiX9Dh32kNwX/P58DcL8dpeh
qg3AhvZCqnCIVLN8Yvz8UgfafnDwK4DeN395rRklxQLKA67rLjQrBkGLoTYyRIcQy4IGIZCSfywC
Dz5hb9I3sEm9QioD4N0Ln/YqaiORv46dl+ySwkzc2r+xYVmAMN+l9/2ovNoO++TvU1uXXwGzb43P
I4G7xSmduiQTofQMQg/tb5acXUv1Ws4nxuvY7hofo6Ht1ylOcTN/n1qgf3Xng7wYx/wNK1Lts0li
8/qAeU9Wd8ZHXTWQUmx75H8/Rmuhihgj2dw5hdjovftc9xH/DbHAv5vOVQDseRm+oiRr6pRgE0Og
5xzSdwOTMsItjKAbrt/iH3DBe90Y8DBXMCErSPrSlvx+NnrHKozmrNKroFO3WwQJQH1BaAu9lPEY
CGmhC0/XI1t6KHqrdOvO2qblZA6K08dKpqA79Dqxby80nudDvCLTTNn2sM73WhxMZ0IoNK2n1Ip4
yemrPLjX0X3mvR+yJj7wiNziISSfSlchwYgmCrNWj3tsc8uSMmhwi585eNWZTpesP1q11F/ggM4m
WeswBOcWae1hHOPActoTqD1sUxX2dY71XbjI6R4NPRXkSfrwnFBCfsbk9FCv9Em/5mqJ35ZETzN4
ntGEtnsBIMKs30nLD1k6WUtP/FhvXaouF5G05FdiwpPzn00gJ1jLEVWDiNC25ZxdSJVG9M3nBEcs
JBm75GYuob6dooNK6t9nXqQ4mm+oBfJg+ueV7dk62AvhMwQtnOBPSEEpogEsy4cdLofqLw2Gl+MJ
LQkQJIF4k/PQEoAz+jbadxh+YbTN/GRA07i/3YcLKZcDwYN2Rkej/JwJAdNCgvigXpnhamCeWG2E
SsgmqTbCepFfTUMIo60xFFTODyb3qpuwBBHF1kYXNBt6p43kM52RaScUClDGPH6NfJCjZ2n3rzDI
WXmxoy49Ome96plji9ofouxh512ExekgRt4nMTV32TCD+fhPW9daXVARweEcuspBw0Se1U5nmeDy
6xICJDQycag7bAjF0zuPsLBjtrStFulb2vdiOGSCPdxvrF5BZdIMsgshcTGkdoB3zk8GyJ9U+rUy
nLu930F9q2y+d2lagicpOwrj6D0WgVPOxq8GLLyd2PfvyJ0gXlzu7omTWEt9scx+6DtxTstxcabp
/mOZ5Mt2rwyFqBxn9jW3ZRkGp6MnIuKw2pEsyLyYBZ2PFuCGTRbrf0RTi36XWP0l1uKKSGaG1vUp
I7xXnFr1TD2gBWxqNUODqnjwYEWQYGo3bETpP152pqQ2sdI1ZGORr20kjGnYYd30H7zar6WcR9/m
CO2kqMXLdE4ib00DxSV9YR5jJnUZdIM0IY6hNJEgQOE2kNlwauHaYnCkrvCrb/R32hjzA3Uat3s2
f74jfzekd/Dz3EGkt9L9UwQCRTEtrltC3zGAoXNn7046hFK9bAIo6cGalbruwA8iP6f3Fm6nzqTG
0bYIlKKAZW7tjaXF4CPReAbFkVISJlzTd5aGfD8kwdOgKeIEh1VzguQPDLwFb8bM2LPtqSWKMUpN
z86Foh5VyNStAz4ffURRh/98xCmZtAnwojQ1sZde7CDSMUsunzemDvF1vLJvWwREUdDTBaGs1mf3
YTglHD8Qn9XBUBl69ZXz93HLdljHJxTcdFSEXiNmUNQAU3AI7lAS6bn9COU7hQKrmr/+xVyvTigu
vSWL1NuanZnVvB+TGTK3rnv93PqeLmh1rGq+XxrMq07ZMt3yOhTeH0/NhjAHwkegg0ArDOt7htyG
SPhWRd0Y5/QL0AVMsov5LPeheB3fSziorWkdgW/x//9oZkZl5Os2XPDusfW0wTGRWaRZIX/uXsiH
iW73QrAyH6py4C+kXJXa9Z/x0DxaztN/Xml1UOm5DVDVqtracksPBBhBQp0FWWDKASJJdJ6sRKNz
IWQ7yBDhhLECWwyT4hwMeNwbDH3aUpMN3zMypdPaRfNDscQKxOHbZ+3sGwvHK1Y+XjpsinYyUgTf
fT1JaYaNdecAVSiKoO0vfx6KzUpeX8jk8B/1OWSVtMPC8DGKrBWKW8PAw5hKEVSoAOMfC3op6pvS
3Je43FvalQSN+vSMvAmVs1pj6aGqmkkTSgFNhfc3k7d1SGabLfzNLSQNzpQndrflTAzgp0o2nQlB
fDp+8J7K1KQ0CpW2wjmaqNE5NMt+Yt5Hsd8+pnw7KuxUZjZF1sO39j3Lw5v8Ml6elbZjAUo+y84h
JFPiZROF2KjyNC6797mf3Py/l7BsjMTwigoQnZlHQ8aWdyUQHLPiGLkmRk9a+ErNVLr23mGal1Mm
oWSUvqaX6M7JpBnecK/hX8qVDpUWMc26aUGFjjgYwqT+Jh75YjbzW52KNdkH7Evv7nCJL5BhvBYs
o7xMTjWVfEHUtHEKzLduv+BPVvehf0N9np+TxBiM6r4LGSSv+qi+loJEZwB2dy6x1IND7qSkhqce
jXQM1zjGzphDd2qwxVb6lq3yoJ/rW+sGDk7oa5hNNVQIc5lKG0N4RMmBnhSHqli2C+pNscjmS8Zd
HGiaw11i5zhwXw+fgAefV/4k2CtUVPWemylxjFGKMNczI7eu0ch4z5JUbOT9MlKtTkXLwS80OcrX
RO5fvxlPTafI0Oy483uUteH3DuQDrlI81CWVdTarmuRKwH7ShPo8qffuLDbLpt5kmvLiO/BG4/eV
u7nA0wdpz+jM/lfJeCw78aqeGX+8xEdgK3eFVMR50xQ8AMpWqFLjTVA2zGzksfGVyhYwvb9GZ/YF
pm3CfsJeX759CK7cPYgP8EmhbExE1sBh++HTbbb1gdhsFHHn/wCFIf3sIbb3XlIBmkLZ2Aun/2/3
rhY7PYmGNWscVj+G9C9bdo5QAlaQ0aKTV9tL7vFfcWKyU/XupAxxuXT/aHrTN4dAzVN743/XxMmN
LbJZLyQKCdUQNbYNDCnwQRJwwBCOkhjYldaGqawst5Lvi594N1J0l7OmDdMv+IqSYfvlpTBmqx+B
/V0UeSvXWK386fmwbyah0+D2qjg5L7fOEArDw2b84ff797ejQszjqFgNB95+yTb3Xz5x31xJr6Xh
gVSmGuXFtTgi9XqCcuLAsMZSKihXw9B6adx+5yNPz8npq4OSwaOT7e6sBWhxJsWflSBAevoqukyg
ogewLiYoSJv0p+8TBJrawCwkZTDz7Ja8ww/Hx4OwoEl8ZKqp/ETdANPivtilbGKia0v2xELazrfD
/dzspmFFubox4IIvk7X8piTDGxV2gKQv2djaLjLYMrIrh3+w09fMoSRIDzA2fzPlzhXzpeTm3K7A
0OKszagrVWIRbAWN+yViQEaqb8G7xr2Mpc5M7dVx5cqGLa+a8z2hHZbbjd+PemN9uOspxGVJB4Sq
Ivhal5WZbWt36eZmagHOAeZmjA6h7JI4bH2b1yfzbcn2pbFfatwdGAWDGGsmU/GY/luaa/PZI+/1
Id9bfgRejnwRHqfj9rJFctlrz2A56uWcDe4Eag3rH/UZZKiRqxnMw/IXdhJyqBIUt3FQOlOLCgLs
9+qccL3siAnuoZSfv8Ybu8W5ruRx7VXsJguDLUfXSis2CvFnIauKRex04KEmNzPB/fmglO10Ho81
f7+z1Jpq7X+hp1wYFbrza749sp2wC5w/q5GXYGsv5TZbbtvOD0gDbGC3LjomUr/RfKF/heaxUp4p
8p5MxxVfErtUmEYChB7VKjdgiwe56pSp7r6IQRCYbAuaAoLaaAmDOjRjnBw02a55KJokjlhiAJ9N
TOTDsitKuJmm81oYFx7gDx26k1WGDBBB2UlCmatPvJELdQXuHKfyZPnqIfKjdd69I1C1AGBvqJ6f
PKWXwQze6uHBOUCqt9Yr2siT6PopJg/DybV8ppJ2nYiZKh0ItqWwxAoxmVs/vzGvne+bxq5mi1vy
AhiqzwytA+YdsSQBYnB2TO6aTwZvpS0mzlZwD2X1AlNrqnyB/EuDP9PA2PH5jr6AuVr7/sPUC7HN
yOrOC5WN4X1rYUHL5T+Wp4aK7i8/UIWqcmU6uzjv8FFjOwI9NmkzpHyp9usvZO0clzJmpyz+50KL
IfS/seEqA8Q6KzKgLYDbskGcayMlfPqzynxjPOvG4fq/xay4pJvwT2SVUz76jsZZQ76b7QDs4T6h
SGV6k+sgTxnAWxWYXQEUCMPs3OS/PjVLXz663FupbewDsRvgqW0w3fbuOpmshQG1nlSNNlYV9nKo
VVfi9rkGCC4TSR30xbiNLa5KO1Qfi9FXZEe5z369Xz5/30lmclhUoq15YZzIVzxv0rACJNKIm9HR
xCk42ryG0rqKdBUQ57bYU0vq4BAq/vQi3d1sqv4dHaW4VxqV5S4AqcvfT1APr7sNcgHJqG07/W6P
90/ExxnccW8PpxY/92NAkHw1BqhhyxYnixZbSGCfvlK9rgDRDLvoin6fZ7JkYGtkfHCf9fPERWKs
VolpeQ6Wf4x9By6g3YuFVQa+XCw+oSH6hCUl1aO7PpruATN3Xk5d7MGHG2NvnZsg0DVoudlB/LWZ
xCHq9CkW5ttpBHhlAnzrl7Kc1x5YUdxSKPKexs/iC1kwK5/F1z+t49Gkkdehy2NOajSIXSEtuN+g
TTXyW117HigbITfw65HcK81c8oqg6IkrbPLhNgF/sanMsbw32FrZ+Ou31iTkFSVJf+NiAxHQOiEN
ZYmLYxpCzWyKe++ceaAAY5EApllFK9oiSpF2y0eeOGnFNAgO+LbclhrdUhcqLsTnTewHz2LK/j2m
I5JtKkfbrLILmdyGzvS7W1jFacz0IF5eZyLWCeYVNrqQeXBT4ETnzgkYduG0qKZU+mUDb9qRQPVq
fDMS7sTQZmC/H5C+Q9y0Z06dINBQVrEmfbV3GyeR3t+TikdHgqxTSDW3Byg+i8fZSkA6lUY3E0HA
84c7U4vDd5saX6C+o9haS/wiFsK+yCExIFKCToty5n6v4S6fACtwdCU1VxBjk1Ov5yUPq0zE2rUX
+O8qSEfC6xWmygNBIexL4WKFb4uaga6Ulpdhjnw2IM4BBqD+R2l9hSiOHQYIJa0jC+PKW9HDl3lH
xNELeEU79IJWtKl0e3Ilf8f021z1le4MIjr1/0UeU2kmr+/Pcy5oUQq5uZpiROogLiOsicQ6uuO7
n9njZ8DMhpKSRA4nwlek6WvjWw8a7rDlGNS7KNErYjg9LESMehRk5JTqExcdzai1vq8ZyyDt2MSe
l3y6NG/PtgBkEF1DAvzAjobDv24nhts5TezOIUsELv4PQKQ+JmiMpnJ2uF05MSuAn0JdM7crysav
uomf9LmQuLnsBCfTgje3aaOx6AVrh1RUNhYn6Uapd3DWBuVwYjFhoRZvpzjuMrI12dHXJj5Ki+dD
bQe0h3O3eykr1wk72eTzJEGCuyx9hIjbq+4TEb6i3zC14SeKeUAmNW9jkN2TaX9WiXdAGaSwxX0A
5ZMPY5k4+X2DdRwe6xJQQ4B+VcAmAZ8S+NosmZj0hWUb4fpbMoCWlJDEOYy3Jyg5EnCks46fmL+0
1qLUuBOhu/NgLlD6n+jkPR7LnL/BGsgmKHWAbnZnz1np5KLdNBWcFUTLF1aTwQ2XXAs0gPKeySpp
LFNxVJ76KTjKb+SUtruk8hBAs1VuoZFc88mNgyqwY7pnEUJxRAy5SLt2iDBg4+NbC5AKuoSSDKeb
8sEtWI9YytO/Y8ejHfZKnpH9LUeGjSPpTqecnEvUE+IHYyEFsgmiFUs/NhqC3OQNmJQolWSSnC4W
hFhlk5reXkkLMUKk5/Pd00fsuEhFwm18PCoZeMwt91lxLNrt456jMYUx+6kJs8bS/McZVOejc3Kt
LCGc+gN/8IlRK3j69jVkBxBKdXrfRl1a9xLyPkR1vsw3VC1R1szcSIOYI1BivVWKSO5LHMrlo8sp
ynpuBzgvh8IBcKsMzbGHq+ZImgkt7/nDnkLLvQ+YAAvba1laz+nfm1B51lg8dRvH/edwWrTtmWRs
+CwzXpuZN3rcR7r3B7UBNzPtaPpXXGLENFNE1e+x8pV4dSDlcbko55KeIFPqPEp9rfpZU+gBXopR
h4clHu8lzcjhzLE4w2i6YVdQoNS0NxNWWxqtpcsru01taXeRYECpgbnmQmFRUWevRRLHiczCTczo
24h4n8Zu0A5lZHooRPzH9mckmeiSIASZdnBr3Pz9VIc9vmBM+2G1xvHztJMEjXvkf3SfEvvTxjkm
469KRp6PRdb+fz40/VFnm8j18uLfCbGnn5ARkXZ21vuYJ/6LJAocUgEFfjPcJMgGImk/UsiO2U5s
B/IsV0GcRE5Qi7KUHDFM7iY27PW7yJwl3AYRc/bHKWB/P5wmDfFpsyHBnsBe1bERHTLtBuebvjFm
l3n2YIh+WEyJMQUaLd5RtRrQWeZUbtIT9573HBNzDjZ+1AOYpltFfFWbTF0MeRMLE/r3ZV2P3B42
mmwpZmVPV6hDD/i1+YINz0Nb9b50HeFY3v1fcerRHn/ormu3lptf9avJu8X+ao7b8spH7lqWYx73
1taFJJIxBhiFq0JA0IJM9qNUoDl/Irmx563hjbP/UDMmFK8E9dDyAwSReHCj30rY85jPGO+/j4AZ
+sI7yUAh9CpjArcIo15Vw0xz1loFehP915UnlbnFJBB8sPbbJ/jo5xOHNeT62F92w9ERLajoAaDB
Kyqw4VOJafh9oQ8AUTdnAU7UO6p1IpDLPsbulP6Exq1bbJ8h3th//tQdxWNq1KnCpeEqK84i/UpC
IfuleJWoFYcIMbBfxdnin8sA1Q9r8YFYCFNMWz2ZQo9R6vBwy1wSor3JVxqmS0CnKjNN4t/NoQ3n
jMwtFiz7SfipBWmbLlNxLIbvgC3cW2YP1rymoBdGjfd77tHvM9rumW5sZFl2IJlK5LhDh/jrehaB
nD+P1xcok1PI3BClvwQy9gydcq5Ne5da9kVLnc20zP+oPEzz99COLDCtqXJ2zL8/c+x14gFJorX4
yaWQi48exrWBjJ9Nfxvu2YwOTeYG0EEO32orxPh+VV/kUl4yyY0+HES1ffb9Zs3+MKmNJO1UT5d1
sZAD4rZ92m+0RH1r7ghvG9g4+Y35m/XGF/4G/CSmbgvqHSGFFfqUkjDLsGlRyZsDtP/BnEP6sdST
G77pT1RtD4u0OOpqTuxfQ0n9foyeC7F5i5daASo14r9bXyoTiP9sjYDY+YAnUbbftqxrOk5yYU+U
qSSEY49QS5NIZmrd+JeXPLWi39FpZueOhePqRSelixcM4LcL3FpOpg2g/M6fsNGV3W/hAnR9eDRl
iRj3MsZTJS6ymBftUiQL/8TqZkcAqake4BIW+8StvELTTiV8tDRjiM+ajw0iW1+J2hhTghJqkwTY
ml2r3ZaA9sKQZVQEaalzWZGMYePshHjwsavpe9NUu0+Dh2obdzC0rGFy0K+3K4MqtDJxdwKGg6Pf
M9hUciQDuvvVEYttxZlm5wvbfBwsfEO4+L+UbcsJotI/W7bI4MdJx8BSpmsTooCkHyuRCnpmE9FA
BdOObW7yCXY4CsVGUyt7f/3s+8cdogM5musXpvsg5uFwFWAmBgo9n6nS2fHX6LydmjcePvo4GWug
wbL1a9ybS/2dwOJfHm0E4yASfuGCvIi9xfRURY7bTWrj/QeDSyCiEzvCPaWY268Z8IGnhKIo9LLV
0Cr0aoZYoDG6WRy5x5zxPPDEtrJn+2wyBMEEbqTHvepbX+hpJ6jZcVvqUaM97S/mB7tYZNiXF8Po
M4WPdN4tdpQwkz8truUdi/Mq8uQx9pIg6fI0dUd8q6/UbjeDq1Pg+ZG+945zKbC++1VVZOITkafz
cY2NvFdgBOcy3AOULi54TE+kUD8vrDcq76FTZlEWzT1PR8GpyMwRNfqzXY/PQSBgt4AjwO/bz8sY
/Yerj5Qk+0Ql3s9ELNhIOxPlqkA7rHchmfpSRJDBgZ7pi7iDrr4RqrV1VVW/kzoE7w5wm7TlXDnJ
DgXOQcIEwWoAf3ox7UgOzDvAk5cCAz0P/+VezCVMBX8vOj75/Iz0td4vdWrHYLJ70M2+B15+/tdC
AhJ+fOnm7X2pkW+eMwP9ARfk9fnrwg+Mw5bDmpjAT/NlSypWp7PGotQUCboTEd8j6DUlj7MdPobW
I1+dp4uF4NFzGXHyzMGRu2EtHpUhlQX+Q50c1WaiKPlBYdaee2KY1dYs9mrVWML/J+HNPH7AxjEv
1lMD/MmEt9ehrsT8XPOWSI45VAMfhoJfSyKItK18XxGUDYj5cdhd9Y/9sG0G5vEUPp8e8ITZiV7l
izd5VzOcCqF3ffoEg/dWfBmLD+f0sUmKr+XFZqZoTPPKyI3mX5FHC7Ceyh1beCE+e2NikjGKBgYi
eyatG1Kjdj/y2KCV66X+RgOWiTDicFNdCXBeGOW+w33up3nZd8HZZmH1UbHeruObcyqnNz1Tjmf9
m3fl6V9Bt+KsouEYylY0AZHwS7Xu2Z96EOAmJ9+DWxkbbcfmeFrY+Bc6uD1hlljQu85bZQk4NmCM
a17us4KmTQ0QByx7JApW4pifM6edX6+wZlr5wGAeJXOzNRqbV4FfMAGbJACMp0ZWNUrbApyVy/WP
JV1Op73ZkYFOrplVvs8f2LrsslcdpMQ1IT0/fXrBo67UipSpy8o9Z4DPI/FwJQWrbFYfYs8VRS6y
V/k3gqh+mbcFKNylGcWBAKf+hOHAuA7/YdVOPqWm5K+pY2O3beT2Qhcki/2XwX6toojQSyBESUlo
uquQMMYmr0fNrbCQrFg+VFMh853EoA00NGDopc7smV4uW0eurFHcFjwGugFYUp0H3P+aXNf7n0U4
RDa/h5EqBzCfg9ftHmabPZvCT0iaosyUIK3sv8XjgFHzDB3WnHNvNVJB6nSCn/3UwaMicPRVXh9w
8p4Ivt+NT3w27/Fav497UYUlCv4A6yj5swA2hA47HbYgNgZyAE9LqahEAH4geFsq+/AMVfj41Iop
g5/6lWX8m+1L78zcoZ/52Opx+MFoh2oFN6WYakRGNskJpte9Og4i8/eLmkRvRSK1qxtW+1MSD8YC
2bOja2y3ckEwWNXxktqSPgtybyYzCrdAEmTTEwCsba1naFU/kc+RokwsxW/Ms60IeatZHhd96uTP
yjYZ6PASUDPmYXkFor6rjJORyCVoTTT03xPRcd0nC9m1jmjI9dkxCEW5XTWWLZkYzhniiXeqYt6+
XyNK63AUx7cRVX2Mojs4a2XV/dj0XpPNSWkr/CIGNGxEtcZcwYywk8Mn0U/BmjMRufLIB/LiG+7b
t6xslOtxfzqOQUOG42+uxkfEwFLk3dlkN3eunEjocilLSQgFNjE7eHj+Z/j5haG78IeZB2TFoypW
2Aqbb7H360wVpJWBolfwySmdTaL7NKXfWSkvyLO4wWtzFVkKzb4NoSLglTvBS1qQoKOMdbaS+q5W
yoUl69Xhy2NyZwVNk5j7T5vd8TsH/GsVczkRlz6ukKghQV7jRm5OUaVDb8boH57wX5YqZO0qqcxN
WNh8GghapxUOfbTqHhKWYJa50SG9vM51BK7AYx96bFOUJ/UMkNg0OvCYKRHvURIQDzWS9QRADZkt
LeEnvLucejxuXbfMi+DdkPZ6xXOad3iclbm7fH70cfogKkdSObT4veBqq1h5L/8+mNcfu4n56qJF
dHti4dXCeO8hAVhJl7558p8KUEPEHav9FeSu4yb8V5oZlyijs5qppsdJ+Y7t9EXuqACICQ63m9UK
YxONsryGnKAfph7TJ6UeBprFMuZ2Ot7QZ7d+sBc2WD1UG7/0F15oRQPZfS2zuxWtUKwCHbfbdl6k
6GKB4hmhwf7BKjgquBfYi/CCo+5WNYkUWV5IRoMGCwrBY6/0Gpd6PHL6tTnPGlscF9VuxgrN17ES
ww12bWAg/5HhW51GIHp5iIuHKPumnON2q3YlEEGVHlc8qpiIzGnbtJSYYhHVMpSrFP2yINMldRFt
Ld6+QFnyez/vnZSUIzX49dSjfOqBwfU0RjAVJyITTCBG9IozxgWWjreLDKvSnEWBpUjP9nIaEQSc
RboE91YjojFK/BOh/XtXEpNi6mf47skhuuBnuFlEZ6YaO+tdQv4vRWciS50f2WKw6RE8bI7Xyslo
DOhBhSncpEW7LLFc4vZIAuIyv4tiIkJezYHZObiu/jD2j77jsmMrTnJc1wfZl3Zy7oB2MlGFRaWG
siDB+1SG9v8Yl+5HBwtyLxEPuUqUDqpAmdHkga2sxDNO9/hx3k9jcQ6iehr3W2NKa1xeOxJdqB78
HhISOFn6pMI8cuh72/f2PP/YFbPOA5r/q3ypARXLhfLPQK25SxUDwgQ8+q8L80iWyyc9MJw2l0Kp
uqHY8jyac4YVFDaLTqJK1PhBFgAGJJHu13Jw2LfR45xn2DWTG1QpKNjxLjCOCJY18/oBOZ/Bc78E
DcLw94h/FNbHh/UQl5BaJGtDGnqxHThIJ0igPVPe3sYhTPE0ym6wdS0us3S+O2e/LwYruAItKpKZ
FBXXpwjA8mQxZoqRL6QXkcfDw4as5qaStewE1+Un/vsGD05BAMd1IhM4SqQAfp4NxVdOxyyXJk+E
J3s52Q0SCBxoy/kh/G6U8fwkNEIT9/gazJyFgI6AfSqsOXxY3Hwf91CKvhN1Zh6Ibsj5SPrHqnc+
5Ibzy+9IZUfrKjLzmOSlR9f3S9DotvRQlsYH4/ZBhSFj8yKbixgWdms7K7MSniOOpvpk32YOw+qC
XqmbUP4FalKWE9qI9YYizIOYis/PLlarZ8fCFYLAfVOKi3jzgeQMYCB4LZnoc5Gg/rP34tsqz8Qs
pPYpB7jLDwLXjSmB9bn8r4cUzJXoW8LR3blHIhDdWnBhgS96wOle/Pzw6K4WgJr7aBVkrD03c6gx
E1h4Ls/Ho9PPds4kkpdsvNMSw6yWzW1iWwnKu0usozX7PeYtH7qoFT8hjMj2jgr/psJPVKh1TOvs
diS2G1dsEekNHSjXK3dyhGhqUwpkcBwCwGGQ1Fsr+CKJDY5inaJcfYmwClRgHIz5gDxMuE567zYi
sIcnLHT5Ifzw0C165wBsf/DQ9mxlXvdK/cdONgTSQ0yOdeNMjrIqyXSjXyQIVt5xjU6uYrdKFakK
QNwnAMjrK2Y/ekm2qO28ys9yneoraCDW9Yr+svj+qAL65IlSTWxUDfKz6FUgsebLsTNFTEhucvNd
Fwxrk/Xh1pKWxoKUvBrvl8e/c3JLJQCQLb0pMn9RP2Z8r1Ss3Ss+jSmqpEIrzyby21YrPbvpGUdt
HgxG9r/2Z8NIdQgzLMaMFHVTxHN0ZNqOa7Ph89RcnVKNymr4L9cSyL78DtAo627ZlmE//5T6FQKH
oFrqM+VAfcQiCq2GN8h4jO7ZIZqDNpLrcjMhMMBiNBFJNG3oKeAYkq8VFdRaU5A0pDKohmNf+FIN
zhNESCKQCDmfa8lgG3Krh6DiV47JpmHfA0tERGuFF1t7sXJ/I31TdzVPmJgfnyGJs2uf4EzS+Owh
SHFEMJ2DBvuDiEveAKmLQWg0b2nsor5Rcia+CoYNjNVhlj941j8mvVbORciMSw4dCzuu2osyAB94
OyK88J0HnbwsD9i+MuD4een92ZCfeTZzrj/5NfBHZi3ylsJOIJ+yPUgWmuKLsO4f1qu4NtXZO36c
py4PZHGE90vkGEp3Tul/m4O/OIhyV+S6YdLHpXkqqFkpI5B+WVOSb4Nphs9dmgWfg05k7d5Vx4wZ
3GZPT4qQMHZvLgPmTYCXZs8HjpZSrr3HwSkZoE+lte90OF1PKsKDOWe3UZ9fMd6WrG+9+VLXc3p1
gtLvyZXcj34VnNrtg5UUs58fAL+fNISRDLvHylYzRPQaIkn9UALqVsiFzUc1nO1b+BrPnV1hitXC
kkRqODMU6xkIIY2eqHihQ6O0f7ALNo2T47OlhvJJz8HT/dHgOaOjmxSfzVvyYMF8EHFFOsMeAW5Z
oUhC6Mo+2FyvN76B2QCFIbFpT4lFFFK+BX42/nBzDiGn9SeFK2MiXfRi1IbHSzxaT4XrUnv2xSkz
ulca1vZ4RlcoAMizB/LVHrAFR7SViPtaY1zHdqI3modUdf8zs8xeEbPevo9Q5xfOS1o5GvToxDGK
1cETSRPls3brgof53fq83Ml7Df8V2WkI26vikwbfKbq6MkzPGldJFgClARjiMzMkSKndxdYbB3Jo
AD543r0UjcisikOfBeQkyWkL+dDibPrIVEvgukmLtdPIsxoT6oftvdTq55JkG7moGlhqN6q5T7WH
Y/k+VOs3qFByUwltIqLNWUXR3K79RRTj3+iMpcf7wKe5BAK/45iLmdLVYQ2HSJD2TsHcz/Jv7Pxa
uB3kFwTbshxR5UubqV1i0QNjPb96KMCz1Rr7rJjUaEsHi6lc4cEVj3jAL5qQwdHwDG43DuS0e94/
fmhSft+aASluVuIwCrSgsfMzhftsw4Tq3fgwjRkIcgKsrrLT3h5ObNt2KsGPAkm17rDAnIb9fNqc
4XH+Blekn8i6W96JEapvVTINDCuiweRfz7Bee1ba94o443fZto9Hss25qK5fX1dCgMPB2W1dzypz
5LdrjQHchLAU55ddnioPlFngAbVKYxhEH3/bUhNnceI4FjlgjvbOggEkuz3jiV0wF1Byu3UOaqps
l1xzsJqgRkwt/v4K7UIMVke0d4p4uCu75AkMwQO6JtDX5YxAqPdCk2gLkz2NKuSI+FiwKtof4kfW
ACxX2mokpmiwmyV2rESkPsNYcxH4pHfJsB4qqtb1/P/u+ScYvLjFIFWz50x/lR18emv6J/Gx4qrL
hbcBXwAg43/Q9tzsoD7Hfc9b3mQg3fyOtneOcNU7AnOm5WcSW8bgUNWvnz/T87Df3+6PPxyaJLOf
TWCtC1AenOiic7tIfP8YQrhOvInVtYRnSw6WJMoaQ1YPvm9oijVRBHun+Q0ET5SiIgiuF2pwt7Rp
zGcaMZ3eD3zii6zkeyu+BEbKFAQR8H1ZdPwuy9HGj4OXypNuPBPFKzp1jAkt8dsITLVaWssQH2Fk
9jtSvZWT5I0v6XyGQLaOHH9/s0BbqOd/Cvc+DgMNQ4FgjAVHB/gW40Mxpk/PDrLjYBkzS0Ep1/Y9
XaROgms2QFIiSGvTUs41jREYooJy+F2YlOMocas2Pywf+tuYUY15W6ePD8JnRIperQkmNH28PdM6
wmfCq7wKaDbf4AwtafVmklbFTlpSoPX9e3G6ualp/NSMOuV80yeNm2phYLkY9jdLuA5IEx6L+vn1
PQh73MXKFLVTaYAuSmE1prvqevHDXKA1Up1OMGEjENDF0CzCyqlHlBsm1u1Ln0o6b5tTgLRLfeMS
e59l9ttPU73fajTeM9qJl1Bq//VA1iUvW4rjvR3BypqOVhvvN4h+7JlLD63bfvbpC4jERglNsVeg
cYgVAL49srYDt4cr9/um5daqc9I42b1j8W3a87s8UyAVChKd/pUKbr17b6LFCG4LvJfo10Th57rF
8AjeEl+88pzHoSgpkL+xm1SmgFbmif0QzN8kDs5zoUf8fGa7xy2LDs6iiyWO1L+5awNesmhwS4/E
YfsXysDXfvjMgsld7daurmOqPhjSXBmw/9C5S/49j9qhW2LXPXVNweCnWhvt/RcM8RCJDI5mDVWx
T7bWze2QVUvFhmaosbH6dbAG8A7DqgNPAdLfeI2yPZHMpuEZ9kvNoRI5ZeczTNHJLxLKjeA9Ka/c
KTLUu8CtiM4MaMrw5rOvQM8AJkEy4WZIf5v4CxnIakvxZQaXb/HiwQsDRQ5KTgEFmGUPuIajN20l
OMQq2xF4wXjdK5rqk5RAGaMZX1LqsogXexx/RfbkHZKcPnG2pxKQb5jgMRHFbx3xkvAJZ+ZsUOMl
UHwl0Te9fvf4eYLFgaoTBOI4RwvNLugW7cs/wLxyGgaWjMtQW0pgs/x9lL0REGzESl9N3enSnNmC
SMOCDHD8pNX/h7A4gfhy+tjf18L+0zuGqvtfuSxWuyzGiJNWk1a3Y+5A8ZAR6t8fS5VNgvKe+C7J
EziDWlASmK9Wb/MJE7yXwVcyJ7AyW03IWRHcycxuqjQFLftLpeUK92L/ZhN5eYZBK5vcSU4aOrwc
gy5ZYZgCE3kyUr8oc7ZrVKyK0ZcL7nt80KypPc65Xona+viuVUng1YCtinahhtBP3tVVJmPaA2Yl
6NS+Ui6Z/a7C36wX529/8jM7uecPL/2Tz1umAyHWTCmRKqE1nykeTfx55ZfZDsqDTTJ0HueRxIJF
GS0C+nYnVjBZBFOxjO1hzoQPPcMKkydn18SjQR4YEcz6rCjEui0qeEmEc2rjOQ6HbIBj5p1N/z0U
0Q+bXS+CNf9+OvxXMUavQ0v2Is1VwhmQC0RySgPgjqBcWAlzbuFYXjOldt9sXE8Fq5rpnFxamCbT
+gmWRmFobhmmIcFluPiHKTzCZ3DtbMCYkV1BH+wSDzGIOcbaQC2FfKkfiCurZwY8/Ubn2igJhRqj
ZL+osKXfllMrUu5YghyXmyvMsJbZ/74XvcaJL+Zjt50m56IGrLmpgUjeoXtXXLGEMh1DeNeOsF+H
cUH39fgQlXoabWpz0CasHkfVuWLSB3fF5pZtZQr+QgJZfQEjr8q0S+3fB0AtNSA/m565PcTcAL/L
4Jr+vNElmYPrOVE3EBGpGC7C/J3Rl679mkrdg08UdRVIoHsqv84dbcBK3fPS60V+1i8uFbUp3RC8
IRzVsAe/14Y4S3jtAq9ndgv6tnkZhyaAahNC2C1J6DCgwvvpsvibzma3exqxfg/gAz7zB463WWnR
M+GfwpMUVtH5W+mLPwK6yXpLQXEqxV+wta0qM7z66hxuXi66TgY5MAlssVnhj1hvlsPPExKT7Ioh
K4vTG3eOtxsXRIeK6sBxlCQTcCyin9PjjAEPoise3DFXK4MuM1H6kR7pbgl5yiHuo1efiiXMtgEf
9Iq223N3BdZf974VzZB5AIVDOaEgyVKhaevtvsho64/W6MW7+EQxvBD6CGIXjDIUDY/go3z8cUUJ
3YMhZTMFTzPg21uH4afZvsYYH5vIUyel7S+mAf18AnCAXOeeX7ey1NnZmPWPIJIuh20DrGId1u0f
SimHj/PePLz4jIcmYEOmRK68TKXXR/Q3olvavSU1NjqIBTyBMzlaT6Vr+GM4CCzlF0KZJKjY4SzW
BGzCLsyWExsQK4mdN6dR5ygvMgDsd+Kknu1iDICBNzug3kkHHJnBiYq68q1vMbGIDYSj86a625EK
Y0Mo+EZquSuBeHxkG+nN1W5G28FtikVJNFmJVXxXY1TSLESOhV3LsKM4at/iIR0T+hFetBHwA65M
X/QCxznSnCnid3RPg46szQ56dFaym9D+u5vXZkb/8tHnHJHD3n6x4mPXA7cg3EudQdPVxJkY9zCf
W9U8vP12ChbQ9B7x6JE6XmHIUywsbnoSbsAwsnj8CZabbIyNTXgYKKblLb+ODcVhJcVwS/kSr05S
GwugO4sC7K4/V3eXrFkvN1/CWkYwNT28RBwsNBCgkqA8PJyamPVwjpNkE0O2rLOjeDqueuQtkmmV
Sje6mEmZ5FC2RN9GgM8g5IZGDLRGLeN6icIpNISyF4BMLpXxY7FeZPryx4o4fyVZZo/opgmYiTCw
3MPqxbhQ1/pg/QyZT6Abqly4ponFnLEmyvvWBZL4JIlUwwWoKi9KMMotegas2DwIII7AAfsJpN2q
oi6u9Pe6otuvA2/P0BKF/5GLrcQw/W7k4QPuO67S/U7aCKiUy+xKOXsNQZWBleal/+syqBgVxy+2
gkZ5VrxzIUG1pnmuwsGGDyCnEhBXQ5m24orC55/wXVV2xVAGNm0hPocQuQyCARzMjOHR+ctVEkk9
dQKPZpjTO7Q3yDrLkixU/ceySjFqwDlwRn17p/aAliJm+uw71JVgudusicVgH4NllOgAEqU/CKEp
uHMmikJA/xnVbnrRLj/cOMehSwpzE81bYZD5OS5pc7V4Sf5VUCAiUrVpUvlISmH3858VuMyWf8Jb
oLLLfNlNmK/rdWGfbsMqNQOwvo8c2c+Ed0yE3X/qkBQPpq/kYk8udmpbxuWAUD8zaq+Y1r8pVR+S
9VvENTUJkp+2U8p24ZgDhwE91FmD1V24Swo7ZhbHUyydQXYstU460nIWZAxqHPF4hDIXAfCUH3+N
/I1BdakYVi2IH5leHRwQ2pXA8qdI99Xh7MZ0TC/S6/BNTRaYDwgjXnz1FW6S6trXlFR49tmSNQs9
oJN2s156TzZ92ZqVzwQTHBTMWj43eh2cnJxvECUR2O1wvMZoG1A/WtQrNE/dbpGAirE46tk0IvlX
GriQHMDs2mzRAx6O9EYvETzkWOURxEDtvnKGsjcP0nmvs10HAdIb+NKCflNuDw67qZEFQya+bejo
78+y+Fu4Xxh1rfnBdQRlTJp8HH5ghjRw48lxtGH9n3650VU7MY5v0vTPYM54e9KymWZah1Lj8TkX
OAS3uhuxRfr7NPnTKPFRIAMiJRP/C+tFNLDbp4k0E5cT+cMjGZxYYKYycqkdFYO9F8TNnlCqDcnB
a8xGckJ/HCE2Hq/Ku+NPu2jczHKtxnasPbNoVn8KWnMO5PjSCkNrNub811McpsY7PKd9DSG1ip0O
1ETNkrxXbOKGSgyYEITnUT2KQUXNMR8w3d4GHEadjWDMRixpcbPi/BSlzqsvwYEWz8QRkm4ScoN7
oD7/eeot/BLKh7Cv6xQH/nd++vsift8y+1U9BeUhiqDNgI+SLKXDIyijdeyjCYwMviPJAXqUmfI2
pv3Y3/ALEucdCmvI99kH4LgrSb3XyfxCYquNhKBRn/bZr5sR0Fll/Sn9PjYSNWdM8uWnG69Xpw40
9P6w5y/w9cnYsdwYXavypFXRLUk6G56OWNDiaoehBBKhbyRq6V0OnegWETUr+fnNRguqfp0dn3fm
K1AEhqfMejj9nzmNm3GxmKGAndvDOezf+iB0yS93uselKqS+hDdzz5UVdhPDp+zexwKMtCqmaP9k
CHuu33kZKULp5xWesxipYoLxiB/BIYYnas7syh4CB8/Ak3EB0oJpGTzMpmxulIJm0ETOwqmGHacj
YGaYCJOspM2mCkchRHB6VYmVvTjMUlQFjc0wzu7nkL0Yzvjdl5reWTZfTeqBtxYkXkEQgp+bgQ1G
za2mzQHWrfxGdy34KTtegmDCJCETS9OEEMWCkLxe+HI+fAdLbRp1IS829PC0n3gq6sTmTJ4rZXlm
hFkVyVHkMiYYMHT3Y+yLbcOSSDiUDiyOtGHpUqbdolBR7PPxSVW1xikrdWlkdY+q7JLWIEyNae87
V6ByG0uakbhg7G672pIBkiSZqST0ap89WJXxghfTFG9dqEubIxeA78L3cwy9Bk7lQCaBDS/JryUR
x712oTc+vWAueLJnIEu6Bsz4QtIxwcCXyF0s0G8nBGFa+EgzGHyXsPIwvUFvGR2kCQK3br39CmNN
b6obq4cdm6DVddncT7OTz/nzW/IY/j/o0uRk3fOl0TKjvlJCMTb7wbpitBOTDxplIaqQZqRI+4ey
UNqGWWHkT+iWiSBADgMaW6GT/EIjRhGvasEarusHcLsLl6EPoRaluf4zh1oChf+kV6fKy+60v3oz
OYu9T1MudMENf2mc8186nrKiZEcc/n5+oCM147H5r06it7M/PZq6fyhOdv2O/800H9L5MydnOeXM
YgPBPsAz967lIG7wZRsQOO6LFg5zOtMucwn0ffP2ONFEV6WR8dX6F61fff+XyRJDsspjZdKxvBB4
6/6X6LIqS7SkCiULyV1obAp/nbYVAKMw/tbvC2pJe5rYKDLVobf+nddRxmYDk+s5+WQPg+yT6Cv3
zHhR4U0WvYqM7M6HPCzJh3Lgiz4P8Gq/UOqNNr3Cq37WnBQKlvh2SZ2kF4taGB5hzWWRaC2cGs7S
/1SYQ3GN3/enWuKgMZOXvZD1DpSB5DhkzfjweZgmks/+VsZiKsZDn3vE3LqA41mdSmCB9XVUwmXO
i0n/zO9UflfiPt0TusnJqWc9FVr6wt3J4CpwigTvd/AyXEKRPySpc1iOPWMRx86RWqCUaDin5ueK
tQMepPftMjv3nteU6UknwqAXC8CyFczAqhSvPmeAU+1VDVqLjiTFgdmHdP3OuGA6L35XsUEMubmP
kTyvevLppNc9CePc8tHvyfct+5iqDXjPFi0LieO01zvyLl+VWYVc2UyeIeSAwhF3FJB7YaYwvRCR
A76xt7A7Nexvry0b5KtlSR7X2105gSlECR7BU6LwCDX4xuGBjjuqGaySBw2cZIeBYTIIGYO4kaPI
3MP6CSZcyffiqHg/AAeuIMMCvUDCLM1AIrXKGwcVxDTKE08XJe+FgEAe9IImEukVmr4aZMQTmBJh
343CwJL6yyX+fGdET9AFM7CaBNitCy0wGBUbZkfxPUfJ5TuIV9DNeVNkvItrDLbLRBJHu7yH4m+P
aHiHLJXfNwmSxLD2xb8xqGiEzFO5wbMrX6b530puGU6WcdzkaaYOVJ24Ui+2wZKl43jFV1ukyY28
CD4Hh46Zb19a2obA+hgLnAUy36QP3HfzX3FbxaKAsP5/phaRNRp3OFRwlwIP1Fr9qiJMIhoPQrzJ
HyGC7nLJJeuT0FRC/y/HAwyBOhDACTIbc4Gwe0fYt3mst6NdlmCh59SAuTUvMJq0tvHOKW77o+Wr
A4eZlUHEtL/zPRbWY1LusszMv7LdHy3NNpZUXdDQSDxq12sXi9TzRG9Fqo+MDme7EATymEcHqTdY
iiyH1bIybjGeWlWGHt3hE20v1kExWTIGXp+RNPuRMJt52ARn0v3DXjkBLOo/hbf9mfEpIXM8+FUv
D7pu2ZIT+KoLlE8yiA6KrsXy5/P6hlfhy4fQy9dKB4gSoj6h7SoLpsRvOwEe17kDYG5EWrZb5EB4
WRafRZua3xMXMhGz8MY3pI/SfwV7IAQRTuA2enkGHJy8cAJkFy91lAt7lWsPqDwHbgAXC539Hv7p
4jNgg7sUiMWrVzDpu6ZQ9zVTatYTb8eGU+BypBHCWCKqfWTLIFHTXPD4EGJopqz5NsiJ5U/lGSy2
8ZhKJ+Qqotv5lY/hDBWgDk4WOF0CbKQ6VqNBe5kRevQ7IxFPictEk2DjM/qauTX5zZTI9PBJZa9U
e/jPnn/ceMDa8irIaR4F5iO9MCSW7k/3slfL8IpSgQrwGLU8kkaqcivT8P8UJRDleVPT1PbjQ8HW
ZY/FqU0CenPSHXIYooF9lcpsjQetIO4GBBvjKLrNWNshELrNcMUKlVipWwTHhihQoa3vKgvVVJSU
TVeEC0QqXBjSt9qkh8UyiTofNRUzB/t0iWoVnMDru93+kk5vkfRZ6qkx0f5McxfbSySH+e1LknwI
tsgDe6jDNOg1JeYzX/i6pcBo07zhZURyRMO9xDx0U3V8zWGE5qxmoGGDYD1hEikzexXdU+LsGTUr
fYfGzLacf1sFq89inizTdZhYPy0AWwZcGWc9EJuJ6VD0IrvMsq3anQ1Af5Jg4ZDQ2orMEUq4h2lO
9Vy8jg9coaCILO4GrSSSk38iwG7lI6X5cnfSTm1kLqU4MNhm9nVYQ078wRw67KUAgHd3EEATWMk1
WuvDYTSGcDSBigxWcKqzhoGul3+cCdBE6z86eP9AHu2wCUgPx1zNe3H40vhnPDCzTPWKHjx1/xkQ
h/vlVA3YcgFWco8KRV7VionTg2TS5teaT5bU7KrbI+i8etrg3uVFQEhpjq3Ew5NhfszhaquMu4aN
r0jTepLwwCdqLHW7km0hrWOIs4SURZHPhkmyKY6XfPSO2oSbcFedPO7DFVoq3gzScYGlqq7tDrRu
YofuKpMfACxKwEmG9vGv9P4b86bJCYip9gIvor44HFQO5JodOJ8TZQ4QHO/OjKlNo59xD/YH/T01
xbxJvq4NqgEAtMQX4QSKhe05RuZa5mTK3Bvma2w+Q6AejX7Mo6CHJc4+E+iir2n36eQR6J9DhYYa
tpysV006XkctDTt7Ysn8Qmv5By/MuZ7KDYmUCmti6qd8wkmj9dk1x9sMXd/byMzWmQMmuD6wB4BH
MV84YQLKYH62P1lxJFGvJtOR9n0xHJbDYCw1eTFykeeVU3ZnRGAnaykbGC8zHrOYfadRkcWk6AlF
A+2/A+M+UiPuwahfVELWBB6GB5pl94OBO895p/aGA8ssES+dqYXLlv2IyQPJDNLL69AzdS4LBzo+
cq2/SSVK9iuPs4qSylo6XTWM7bJ/BBMb42Y6N92tp1n7qYqFW8BE5C7vltIXM2VZO64ktQMMkbG9
hYSgMeFS2zU9E1mGNYOPi0RI9GzEeFQ/ONgrJ/9gfhC0hfoXR8NSP3LCE1QP3WwlIDItkeLpg/Ht
rF11Z2oR+xGntqh3N99o2hjviLkpZUnSwjQ84Z/Jnj28VtTB+1+oaVdYG2J3UOV6FDdZHcmJmw5J
XVb+XCkrOwbKvWw+wKJWxVPmqm0Q87wewMcelmhA0N0a4UwzG2BFCFdh+9cCC+g/vd1MpW88GH2k
Z+Ae1Cd+ij0B0ilD2KPosrKW9x+bw3Ql5c+L9WZq4HiBgnbqzlHRs4Msg3rmzyvrcWLcoiRpSb7S
NSMSf0d9YvELsmxxruCVHzn1L3aViYMUOEtrIZD79gm3rMZiPoWO22unK8G6I0STasxG/1rL3hsJ
ftFCvak/5OhzrdsRbUsWhAlD2UhlKY445QsUbJwfYavaoxSPagHzhucZaN1u7W68Ey0i2aIZptMP
aMT+8MBBG7YAZenoXL74PfzxNvTw5lOVWFfIVEqtNFQ/RBB5rTRx6gHMF+4XYsUmuqWRuR1fYl8y
hX44D68WnYjYhTKpOYaqT1yCoNo31firgFPcyrXD0BzYNqMqUZnpq4epCfXsL8mzDkwdDyzes5+d
Q6Bu/g2JsNifLJVHDOO1OHbeFJ/ryLFEejliLOp6Fzp5oDsNd2ptkuVHaFKIPR0ziAe7Bkr8mxRT
sd8P7y/jzF3qCGr4ul2uKaRL/1MxwO8n8ToN3J/VvwP2gyLmja2TZOkkzuyKlUlgFT5FW+HgqwqO
ZSlYOKiw2sdMxHkxIxUE7CKHHSXR9ekqe+ifEwrDkcCZRNuVB1ONX/wxull2LTtMqmc+BdW35MQc
kaiMvtCp/7X/A4STL2N2Yi4ktaaKCqM+MtLd5DWY0U5W9Ss9V0Hp0sYWNURnEtamzd67UISLK0iW
T+TNgYBzyFl+3cac1pU34zRR+FGCAiI7nwSCg3sUtNpcJBvgA7Yhe96q5/gCp4i+nBZJY6pxsLSi
pgqeG66T/I8OYUtRdI3JfZO7aJngjFKXoGm0EM5yXPpeB3opHtnnaKWmr2K6hwgPln7ke2z5JhRm
bJczQER0iAwz3fDwjSWKbv4LpNpuJ4elxBJLtohm0PiJsgdJ3UWN2RWZn+J5kpWXvt6oMjD7EvB1
Q9B6f/a9TJfG3dMMraFLFqGgz3rzijvvVq2HaKG1Wq3By8EKW4mAtu4vGBPrKYbeG9x4XCuPUgbg
7NNAca5fb7eNfwR+bNnAa9/uM2z8FNBh7l925R+dqsR8Hb9CIJBtA1kgMwZ/HY01nSkTzI+XOu0h
fKMvqFi8F9RUfKCF2Mebp+qkNZqtlJ+WvsHZJOP/rE24xt9yNTKDD96CMOeDw2qQF6tH0Vxm3qTF
7IPZH9XvaXsr8lPWMzUe842CfSi5sYNIYXONJBsOu4jsVkbhmdgF3LwNGgA95fby1GtvvglDzU6I
pm0w5RkMq4pht2Q06oG5gMU6+/hVRxdEZNeo0RQYRJajEjaQ/UKWAwE08TujuUweknuOQV6OencJ
1D1wY3uYDBcBqstg54LWO0+HdTmve9A2NHFu2QORh2TvGCvhumxzYClyaFVJRSMGwli3mc+EzlZD
sEkjJMdAHvUsSxCxQZsll5yD88ATa4VBiBnJ49RZghOmdPrxz3S+gROQ650Gn86EgxHPEaBXzX1o
A758Ctdm0p4n4Ga4Ngos45Z41x4M19N8FJuTqNrN5JPu6hYPyjett5a2rAYFeVM2rWZ3ex+bwQEZ
9sOlN7s1DTQRCSYl7pgOfxv28foyTPmv9Pvp8CeJE7ZpxgVxjDmK0skKTc/IVQ5qC4n/reGsoooE
d6uwBGBqvmI66acYvXHg0iAqpsrPJyqrgp08XZl1zuNMWNXfR0dVug3V8R9DC04XA77CNkiVSy7W
fAibA23h5O9cci5J08WOI03k62yFtEljK5E1vRFjdJUfkugzdXVbFtx9XzpGk/qXq6gKmEnVqxOr
Rh+s5zNRPX5oDrpo7rx1EEKevzbI3bFD1w6fvDDliHJA4j336ZD73hskpRHeV58EYvJ4B5ga4n9U
4ihERI0fMkdwV0gz9k/k2xdJEpOdKjd07P/yfP0cqjayGSK3nF+W96Qh5ZuOrTodOxt4nA+NtJUx
hYvbziMO2S5CaCfZ2svrHFYjdz5JEs1NWF49iDUG3lSAF2bj0kltwQbA2HCh4Aq8WSNhFk03eSCR
skhJY1t96t2eMidP0DA3Ahc3n8SqRWw5aoohK3oKlzzJTTzWLNZjAYf4HHsqDjww3QRxfbhLvoOk
V2TzdFYuGfCcetQWc0ugdwsR+8Kuht9iA7zm6kwQMAvLiU8bnIIAL9lLbQSb44vdbHWU8q1FKqFq
8yJBYeZj8D06DDVMkB8G29vw2Fetp0zmLHoNiSfyf0iP6Ntz8eyJs1JcP6RzSD1zG+5r1SZ7rmKU
srqKgxItcgfGl+V+wK/0sCRkh2i01kSnlg/EQWYoD0/K5OflK/r89u6o+gnqh0JOezyqGlG2gKlM
K8TjCgY2jJtdL3twSZF4Qt9kNN4df5qRT4JzvPSWyoiThsPqJOenzlYgzO8QG9faB1vEK1sfCvaF
jILo7XL8I81p0nIa2uB2A1XzjWALCTx45XgbepYTEMF7FrX/6RDq28WOc7MHnqSSu+DyFr27q5h2
CiH+CFK9Ecmkq6fVdGRWxVUUVc+Lmj0YUbYAHmmMBwMFP1Vt2nZ1B5RYZGcMgHx+RWeK8FdaNWPs
XagNxSs/EuYvMrfGbDXIQaJpLHlsxmqUOOlmjnxJnFXlpye/X26my1A0g/+VEc1ePBY7YK3nkgxO
UcZgaSWPmMIubDMBP3w5FRr+wvGiVTyBH6yADqcwLPImqoQI843rNfJQoDAUEhNFLg16E5x0DRYo
lH1tvYtURmxBYrdY2o7TFVJ80r1cbJA9Eex08irCX0yyvXNXDXDopCMijNnrMGixDbdPB4NzN43A
TZh/3zyUfromrJxp27CFtInLJ4qf41TAwVMYvP/7yUd/1JkurkQk++w0yVA3Sw1zXOzS8E345QaO
Ky3+zglLpkH4jdgTKv4AKAKCXHIaQt9pxEzYFJor/aM+E7xnot3X55uOGC8fIv9AjHYzDPYqE/OQ
aTw55HBKTLnhVvUUHGorE8oDkUHSjotpZQju47FuMW1GPjSke9Hrwfo7nNu0PaepFI/8GqBtCKUY
h6OjwFyVw8sqFwe2FMoJ85Oe7edyVaOjTyyeh8BXwpcHRJQ+R1HSEGlTJy9UUrC3T/IrTejwjaqe
brSqrD5RsYe+yXLUpq5STTY4bMv7y4zgYpH3NDUSKTGBn7Cp1JOmOaBIuSkcXSNrCgWN0CpxuP91
bjyLbTbZ0NORkSv9lOWUCR9hTiFghELywAiAtRlC95IvVPE92MiXn7orHxrPvoZLCcz9YJu3eNc/
tlGh9pcVeIE6Yov87VvYjazL/v9lihcGf11BvtzIGktGpXSxBjwLgOzu/kwUxKE/Xe5CVGocuikw
YLp4uPaOQhqI9IstlqU3kgGIWBmVqe5x96Y4s0Iv4NnjamhwH213Oeai5N1bWO6xbcy3Wfiy/orf
/6OkOzTWn/othu/tAT4CzT5DrOMADf0NKXPPiTfMi030K+JfGGXXZGlu3cCV7dETDxw0rvajn7DE
dmOPZoxfL/9EbT5EJJSwvbb1fC5Alyg9LameDakQsD4uxUZ+QM7OcZu6KuukX0Adcf5tKr3h1DQG
ufsp+nH+MphkGRlT/1R7emPzUkTF3w3geiZ2crD/qAmYskK72O403SoUFVHTygbdvhfz7ZkhvX7N
YRrHiuIMwgp0kF5KlEy3PU81Nzi7ws14kgFqH9t0FhUwxKMEIlbx7MhqnSUqhUXT3qrqGdgJtHdo
tqyaPM1zSNhlrYJrORuMhiQRAjdtEa0SiEeGMeuKrObqlZDwHJdwDQVI6XOhOPlblo/Ef3PdnYoS
VlHTnBQEXIGVdpDtWFxtxpUUg68Rz5b5uqc6BFt9dHnu5jpvLaEjjc9VoHRnGHjSuydUgLaaUPFk
/pVooAyVrY4++4s3Y38OO1phpe8XtWc9BcPTIAZtvUTA9LiDup+MlvywQ8ftJotKP4I/LY/v6qzU
HV2+j1AD90xvtPWUZclZW5lMDzKqQ7lacFudt1IDjK9V8tE+Bp5c3FSy3YlAv/QcTd4zMgTByAXm
mOJo3L63olJsbjR+idFg5t+HJyf0zO0xbA2foJZgrd8JgazstoiO/+J2F4SPZGArFvDOLlQNjROK
0PcT39HF+JiBAx80Qife0VabDPGBu6Azy4MyDGxV9ZVDRsMpERLS19AcKVHMOKMu4TvXyGm63j0L
26rpW+QjUI3KjUwhEpkh2Iy3qZvnCbc4zmlyoiJPHDYaD1ViYmK1RVH7f1y0zR8+AxnIw/FdJ/h2
ZpNrtaAKiOfgRuZwimwxoxhVeVm5PMEsYB7R9/zPPcpXAwp50oDYzu+ZaODgesbfTOYziIDHIoH1
LaXq/rxUbvnpZ0o19zB7FQo8FFrZN8X86jsSMgkak5y72EZz92xATSYBzI9cDtzNR3WjRR8R7AAu
1pz0SXpGUoSJufwsLHGRD9/CQZ5A53cGmgLNHa1kN5f76659cqi55K5v2EYYJ3JnngO3maZSWLKT
5D4V7NzCr/HxYdhDDKMlKfKCa/ZkhmhrS4+9YGCOolKgHRaNJEJGHA7SGw8OxXR9OQ8kk5lLgD8B
MHHkCKfnE3HhRSFTX5LNHy2M4n1TCRwVWZMJSOReYUqWFAAMCZ8EY296cd16n6kpwbLQGw3/VMnf
IAxPf+MQVf0YedpkjE/Zd38SWsZ9toIXHBmot0y+3fjN1gWo/Ep0TxLXerwD6aJksP5FkvTnA0UZ
ipRuTwp/V7amTJ86fmHklqjiocY8i2s0HyZjLdv8Gt6gyLU0bnwsUKIxEoaq8XmQLAgJqdMZu7D0
sPnS/rdLOS7hfdJc74bZD4umZW2qe/h5HzHdS0KiwfsuoscKJfyyn9M/y8gHivvhNc1twIFPqnaR
+7rb0IJ4/Y99ZGMTLAcZLSw+WJ3bYGQ9wKHMsI8HhsQ829/AmX2Cx15HGAcBwYp5HWHZV4QjZPmF
edFtw2L6u+1WfHnFTSxd8NNC2IJvQCVG3sollhLbwVK/vW1ozgrCQZGVO4znFQNS0KtTEMRP0v+w
WvGbIJjD80z1cMEsm9gLbB1z26kBFOZIh8LD7sdt4xsLP72nf8Cv9WmXIpQczvIJVaBYPus9uTry
k7cOpJznCCt48FfqPdmkScnhpwJmidtQ7jvmGqZHG4eWpPQVB2Ptfq8H39gFpQ48rz4UK1QMmzzD
Mwv3fmKcnS0ZUuv2fJokbe6mlql7tDp4tRO9Em8oGt2CAkZ6wJOH5lItbw9Rbiws9/IR0PSym4Uu
TqTXcJgEgWW9NUjcWH+nz/aBz5Ia5g5mFg3kgDM8jc+U9JVoBQiw+KMWa5WqEGvsdEviURZFo/pc
h2avR03ymNc3Qxbkp/mIP8Zx+KeZ8LjcMGaChxR4zn+W4AGxY9HNYxN2ej7PcsxAg5BMlKtNKfTd
dn4wCVynYlAhqSv+ziHpRknz4mY2f+j6WolhLETZWJccVY2sW9/hJI4bAgFTIYW7sBWCDP0hFZcN
scMmZjq5bA7ePlLTPmb5pzC+1tKB2n0txk2wIHgPYgVjBjldwuxRWaQasJJTUdfdYF07F05YmoVR
xnSq8U7O63Rg+qf05LUdMCdAXlaTGGNEBt1k0zqc7dB935vd4X4ZPiH4R8IGnXawkWQoPhKOyItz
0NJ+3Pk0G1suLZNR10PHTnqvOSTBsUOZ+CvJCYYpg3mgpBnPFtW0zKEKcZtcPHbB0wLoBkNYwmpX
8CcEcNzokg+mrj8rSdv+oO9LUcBbD0/rNpCPZxrKhOuVQWxLQcMbIcpm35chuY4qjCcZS0AurmaV
EAa6UdaMNtGSspYQMB/nu89MGH1RsK2sosqsCuLpLf3tq6ZVQnqhRt+UQQ8lmDkUVVC0IQinICt0
jAY5dRV+NXPU+tAAuaVvXJkaCY0f0snSKdfsSophVXpi4TjuAvdOjyHUtAzrOU+B257CRsFI7LcC
op961bs/Vbo/suHD5EKaR2TGywgAzOEaONh+dq9BMHxwp4GQalCB1KlEEyqiHFVr1N7AOWhcqC2p
/IuOEbtBcQf3ZOXn38k+sO7kjLpNgpwHJeXg4r7oT2BhAElnjARFYnZqdRf2SnPTSPXGobWnzdDr
nJu1Xlhw85Or+7+5+m4yoROj12AggrHFipGelLNM+/P3P9c7oncPnpbc0SOAIN7GrdjngrR4nro8
VwG0LJs4twCxnyqkJhPypaCOwk51+Ov7QIkHPcnWVjPq3hj1dbD/mwnaxkAQty396ZOpMHaT/3yw
LF/khgC2q2tvKpxfi3O9osOoMdaweYnZUyN+0Xwre7oJ9pPSR91LFq4ZVTMoQB9MtkMPja1FiHqL
ZDsVOLDX0iGXbHLwgIFj4cg4GNOuqVrNepAEtp5txxrqD3HgmWw5Xyi7Xd9pEMTAkKyDus6caSNF
cD/+R9uSHfLOMgSDoqWlAOeem/cdDnMCYJ+2/AXrZfJp7VxDMhCQ5wbgIUP0BA3G7dISsgDBmU3q
LoVo1kNfR+6LDQb/6a2WyO8qf6j7XjaAmMs+mxXJXvPFk+LLJ3GHumr9axvZq3J2GtCpbe1vJTgF
8RoByD9DazqaATMKV82FUQuLxvb25zBm5OvOQggg0oyntPxdWWfgU/uCiw8ZaM2ewPvuoFCWRLFd
DBbC5SiKDXDvFuLrjqKf6KRsVesmU6muC70PRBdntfb1EUl23L1y5EaGqQ3yevBvUHoQCBJ4V1bz
AjKs5nrTeuZzH+HNzjt5Lj+xxWvGBBQHbV5nzqg0MN8A4nxINM+GRgQloyeiuG7g4rqrGc2n9bcQ
RDBE8OKvF2wCtcs1IvPXB7ZVJQGid+sOQNx7FncCxWyOvCByeeLeT3I3DCu4nrLoTjFewk7v8/fn
bHgWP66TABbcYBrl+PK5janWVr9xVayLIHiIvYjmxLFzymUfpypZDJyS1aUHtxH3nT2Ff2b4f/dD
JySWV/jfP7r6c5C3Et7iBKyzC45R5QY0oB8qG9HCxTKnC+6TeLj2/jdJS2RaW7LWOkAJmQtr6KBK
FBsoC0GjGPwaDlUjhoYubNDbviuMqn3Ow94pfTtAgp3Ab4SIJxu7pwV7W+CM1sJBAhlj4ekeLFnv
YBR0010bpib8FnPEWa/F175a9NcgcSuGvupDuiP+fx9JKy2df5wS+6c76f5rvJZEHzDR4nNGu/55
A7GPrLqZn/cbsVd8A7C+WKLQXK/2ZGbyjJwSwLWhGUpi7HnpKkFXDY7IVMrYDdWxmtz8NOyDptNW
YRMIHaWuYwYSqyJYIXsXJmobgmO6UFJ3VgB8PzpidH+hiNXuJm0B/MlrmNIlB48v8ufN7lN+pn2p
TFyC3PXRU/Rwxkb5xoy+wKKgFYQ06zY22l8WNlIQ+QTPdgfUG1Y2C+P5okdZf6OCONcAsuD4z1lx
+PD2I946kXFJr2xicS4AxTLml4XVYzqrgtdKrhVsu5Is57oQXyWG+I42PsvbiC/5NBooguW7wKDs
XSUHQiya5jhcuTK/hRQzQ2a9vQCL/+si1iqyI7caPBo9LjYIBO89Qpq4akeoKLrPqc6DOv3tPBOC
N/KERqB9WLdi6epUC0yHmWHcWPR79mFPE22NmXjFnciIOhHtza/ILpGn2s/gpeYNE4YPn7VBizkm
+RzrUKQxoQTMGeuLlCtST1vSxmuqLErVdfVcdFdv5XhT1b9OWjical6Ar8zks4jeGAyQlNQ2hU5x
oy4g8EM1dV0SQB+Igbp98qEk99fLO1zaawOh2Cs1DUIcMO+niLr7toI+kCAy2u+xgvOFv5Y4Y6H+
MMOML2Nuk0YLdXt+YOjgM7Rtkn5m/yoY1K+GIXmCV7AqB2ayXiS+5AIjJBP8dJx4MOorgwZLB+VW
MSHadZiTxj9Aw/dtVeNKW4pkqL8CtGT+uHm0az58dmaM+vE3ydfI15/lJdGJ+1/fbslvdlCB3TdX
62hBkMMq5DJtIoSI1CMEJFHf4OaWxwj0iG1c6wnEfCMIj8m0J/85HEmlt71Ss4ZMEk8RZNm480z+
ywyzykjjqvzbmfq9qIdipTHva1Ddas9s+7p+lWO0qJSIWBHiNtSzvXKufdnMaCzb4AAfaVbeQW12
FKrV9/Kh5YaUuF7JB3msfftNWW6FKque//2cJW+dy191kQJCOVxvAhNLDVovt6M/px7sq6GVhFTA
h37shGnTz6kBrycqCwwoaV8alTCcRJuW8v49D1gIXt+q6FUfF4BdNoPFWdO0nq8Y9B5KejmDTJ4g
XPWM+ieITSE5eSIY7YOq5+vd6kWCNQqiChWm8SH7tlW/fIrMGageEHni8R6IfwqsFx9V5EiO+xFI
I93yU4lqAzXOf69QQMYgDcUMp8fnvizPT/pIvJq5baXeYolOT34fJbeAjL6sLda3vyds6presdnE
LyNoLLu252CZDrmWEDPOQOg4GA5DxbBQjgTB4ls6V6JkHD20qa9uoAJHSZiM+5PXUvA/iMS03flZ
S243/hkAP70WXpKxN+dXmR3tJyfrwfkW86AOIiKud3imUMWaHB6+ttqpDkJLB8W+Pbcw0NMOzm3n
bzlKMexefbm1vmt90o9DbaYZV4WWAa9dnkX4rDyZBgW4zXaYQ39yNOt73butWmDSxMnjZ1Z+waDb
vAJi41ms/efEsDPOfVIdd5VwwBMqDgV00KdmrZH7j2Smdsh71GBgWQuLOM4QsEiZOxSELqIYB88P
Qlu0NWyX4cOVzuw7TCKt2TsC0JvdxwA/kE+jYGe2iFQduqdIIJCKkCXw7XyUNTUgPKyEa5Hi9KCW
z5jcfThETjJXkoLPNPjBBJM7L7x9hl8LwVWmO2GWM1h3/cAn3wYHC1IJ9NKDAUOXKvSdz2Yx/Yjh
9NPh1wLzNp7dHGqTqumKmanMElbAzeIInmS+tWWw/xzLSPAL3ApB0rjauBfgEhNisNBCnz4MOAG6
pY10Urcp7xCDzt7bYY3gWw36GgcYnQKF6hoEYpLQ6NflJiMW10OPXonNt2MaOP0rqRLjfE5aSTNG
8QhsVXhz2o+8obAwFNHjpJea4KVNTvF5SJ9QUzqBT8hlg2mc3bX9uIRmVCi88h6dEl1PGj88Zag2
GkzMxMTOR2CKl2Q7RzOG5XLxtDHJ/VCiEzTKCU62UuI8bjpmn/dUUE9TfJeR8MHPDN4xqkxLc2oD
hS6QtyDLajSGnhst5N3WP/5MgzlP1Ipv36uZm2ZBrAgNtRZNF6MunwGu3V3cENHK0Q04+xx+d3T7
G2wEeks7n3Vk0Gu9UYT0j8MfHdHEAKBHZmNrFZ6yKEsqND3Nw4u7zMY1f815SPB5+kBBRAGQFd9U
8Twxa+NeMb0Sfjp/Bmh9oNvG7dMG2VwXGI4PMkhwmxoezzNQsKUbKI5b5aUuhQU1ryNLOanIXod6
OFDDy/w/ED2mUpE7n78h2w20v4sMat+FR9hl/MjQowkmjhulRg/jq4e5yWfj56H1VxpSWkhULcbr
7pGgnkcO17GhY9lwA0t0D6v2BELwPrxd9NbseEDsmdcMwn4wcfeuDPv/zd6NKy12q52yswRVtkgJ
7oBFYPZN9rocJTBbnvszZh2ILLcZQ4oNpD81YjTaG5ExvLVe6rTusWfANSZhKb7Ndu8QeMKwdoa3
cZEUYsC2ebgR0JE8nE+fpmMm36AhHP5aAU3tVQLSI7gdHlxs+SsBDsoZf9IRzbqJL0UANH0NSH5U
J3TS1IEJeG1LNeCI9uMlFj3a2eGHMoSDfZUOE1AL9QrI993PXYYLl3/IrAmMwWxmwXTq5TghwyiS
A4xd7l10uKHPyuQoXRwEiV/KFzpX72xpHLjNDAh20ejQVvWuJfaoZ7gjrqs1XktW+8MdHKG/cGpK
1WtxGXxsNxn4rA4LSvg6a0jxkc4EuCFEF0vBitxldr4eUoBPa7SiZLGMF3dVupp3ZAzB6mBZggV9
5cLm/oT+MelU2djzGOQ3XPUanl11+Trkfl5DSFxgdTOJ/KdZT7ox71HmRf/GhzZ/w2LFjslwPG2k
4b64EqYk22XLX+4I1FY+Xn23bGH7cTc+alEx4WAzx/HOCDJVe5kvq3aBQMusz6oBX9q7haX+NlHD
bA3sPlmoSjGqeWW0JzfuPfROJI4pQLsm19ke6iUOEC3mTEbC3QoIGqnv9WF3DD7ce8rDs4kMRjtH
TrbvcMmPfUSFF+pA3KMG5ij6qDNlnFYUzYKGYzCcquvFvCRSt9wdPQewxNwaP/jJbxrMOGlVEf3R
tKCsKRYLh1CNcm5exqL+e3nbwR/x2j/rXeCNPwDxsWSYayESRHicizvkehffXUpxSXLUldTkVMgN
r6pRmW4ZtTJzOYsvxcbALaYo8H6HagYkqYfoRwFbG0d2dm50Dten9q1tIWR+7ThR2U+hXFr7H3EW
e0jNVOyECoZ4ZjHSok3/UE5LjavXcq7BVsXOl35oEoh4vVngEUPeI932hgD/A4M/4NerXDV4mS8R
pY7YeOEdaT5R26OeYMzDvoWI8Vj9p9Yx+vEWrcx3J9AW4VMIWC4gx5MffKXVsSpRD/1/+fvLroc+
8SG3zIu4QBAtLRNAv05pSgzs1xYq2F9gr36bMlLYYXWjtyybq0ONU3MKvaCx5P8G0eO+RZ9+Vnc6
+YCQ364bZfdS7gnNEJ4+XAIkbiRAs0AyYPjH9ad/pX/zB4ijdvYBoSuJet+d64jSEohrFqyoRBib
CuDCSoFTTkJEO2nIbfR2vDIxGWevBP0Ync+5mby0XdgEEObz/qai5FENc3ERjY4E8p9towxpiiGJ
z//nyoaOypL0rsE/8+GWoUp8hFh30fGdl9MuV5Xz7dcVP2hSO4HE89OI0KWjiUc59Jzygga64zXY
yDeM0hz5b1w9mKFdMbiw7APMaYU97icimwNCOXq+NarFB8XyfNrqfwvDF0axRMhkSap3DW4+BdCH
13k98+jq+j4E69hsHeOjrh3pHvtkbXfaxg5e6FJfahApgpMFdhL3ryd0rkVXT0xrG0tbUxdZzKw9
ry+8cgc7T7prfm/nSA9nC8l2DMXi9Qhr2r+DpGm/ZsaXJBQFYQBLm986IGgBQ2Ou8fC842TFE73K
IX2oF44mugQRtjkKnIqAhBKnbJXLsS08FKJeyV+yz1Us/Qj8Dfxu+ghF/bAQmNp8iOzLQcciwGDM
3ZEU2M0sNdXID9AaLEF9l7WUOIR1wzEvqwlFmd7X8hSm/rDhiWT6+RZxP5zBOb02Gm+IczL0KVKa
VTy5L0M9BJEqbwdOII/8IBzYy9xHaBR4/U+CWdyM+GUCbZq15JrxJpN0RycldvNiBC749SbK7x6O
x2Zy9tB4Gyl3RmgORK+HVFCp0Wb41i1k4bt/QutOHR5ptIQNfooAWG7dS/N1ugEiwGgCtsDRZo1H
VTpfpTHgqF+RGVMM7YyEhvMEYYVBk1et8ceCo3nnKbyaxtBo9rKCBLJqZCxHuNrLYykpakfhzb67
7wJ7x/xhRJzfVB36tUIQboJUVqom8cRYjXzbpw/GwpJEd0+NBXOkhsXatEaFdCPkVKlnOMPDe8hU
AoALTRSOQm1Uep5GdsQDMrO7VHSDIlCSqrTKxABB52j1iEEEd63RkvyRNYfEQBE23i6pMwNUAcb2
p4PWmGYkqsvuuHIa/FFupjmDBnRJ5dD/YUnqKg8fKtG2ZFU2F7O57vftU6cX9fbZ+x0yDJWudy35
aOYzzCGWGUUK5lVddx+vou/togGAm/iOyzEywp65fQun/Px7Y49NRYnthTl/t2G30pFMNU4VdiTP
pzOLjHE57WHc5nKqNa9QLsK8TXWY4TppvX6CZ8EZowRW1QTQ7mCOy8z9SRrpZrROqSa/phcBcstB
Q5/zsYMHVQH6dppGGaldqE/c6NUEcpBOwBYKbex1+3ZMO03vkLXJwhLfpVj+6tiek8sjq4HoV/px
FK23joXmFmq/Fw0THcrX0B/vdaJ2SaAiznGwm32Hj/+hGIms1QpWR0W/j/raQeNzGR0Xwtxrhbsy
Mt21xANAUt5znTwrYuiw1mnzRVeXWaNOCB4+fMp+DzxTUcjg0Esyj8ZTFlHzv94fQNdl8DvtNvgZ
4YxMWWW2Jh7zm//9amuoSAZIPYvoSxV3LJnb7fikitFxlrXR0P9gIkEwtEuoB0bHqnfWCFmxRPNW
ot5fGYsZeS8SO866im1RGO4cOZ4ESIBEbkDuR7zeWIjG8NxM2CEReOk5/pNoqGGBaJG8rE7hyWUt
RmpJ69DgCDDezSQeVPROxkBwwcxUmwqsJtf9UxNduFVHnIlqvMt9p03BipNXR3iORZEz/xyZX35L
GN1s95Bf4Ok5PZCUFyZrrQgjyN96vKfz49+UkJLBIPN9x6E2q3+4c+B+Mlw5X8K2x29fEYzNETKy
q13q5vm9NXycJo4LZysmAP3PmUfMHqqHTonaVg0svt9JSamMWHX4KdOc1XGR2hWojsm/sb0lDHid
cv71u0J8dNzMDKNQJmfv/30JyXmRD+Ft09fAVgBqIO5PwvmvIrEK3uwR22JXQTFZXcAOkgfcXckN
Nm3cX096bldAguT5FYt1fJ8LPgE9JlJSqyOM7McqEAvv9dzkokVf5czcyPxfX+BxYXx7aEOcwYO+
JhaDxUKVipDIPNrrCepDkMwsVXIJ9B5OQyAtlWi2WqWC2eG+vhl/fq29mjTpWi8Pdv2WwY6HOIeR
ll0uQ3UiYlRpFR3jLCMwlQMGW2HzfyfdpSQ6VZt6JTm6cd5/u0u+zLh7o/0dguAmOcMVXg2UwGnB
cLAG2nrg0znRNK+2cfZh7RGQbei00dUFfu/UNjM6D1zPLZT0EXno7wD6y2mPMNkKFyVuYPNka4LO
eiTBF8luZG7w66Wek3pL8wgcTQz1qU/O3wmSBQhtTgJbVF3oSXYheHnVge4eklW9n/mvKhPE1JHY
q1vZJG2DPAeu3Zuf+pyskYs1lURuD0o28U6wyL6RYZtxx/7dOfRyHfzcTQYv+IR07Mg+gqA7DmGn
Sl5R0K/lnpEekHm8az9fSchQZRiKqtS8Wi3aonlR/+qMbrigJhe9gnEz/cWfJWIy3OqhHN6J+VSA
+G8AViI/5QLNPavgUEZCnm/J9h5gV1uLt7wa489HEWRlS+PUKkYG4aeOtuj/GNnv8tI+jARDcXKi
F716uA7OLLd+X1Hi4hBDub6Ah4AGkdO0pxj2q4v5wpSNIJfqx1JeP9+6fmKzdqRJOqMAPjiWmzHz
kFr8uVtEE3xOnv38Tuk/nhY9Gu4+urnyIHqC/YtCsSxprBi2FOIQ5RxCcieVbA6PXhSqnPPp+KDW
eSiB8wkO5NvcHfoj+FAHmJ6/akwPXK5hUMjL8mOBl98Pd4blK9q+zDMho8FrX0qOJ8/IzP3t1egz
rukONH+2s/hXlVeHT2DBcI3Flj4wa48yZBCAR6F44aZJp4C4H66ZoSFXTcJUKCTQdn9Kb1ZQTxEn
0RUddiCPZNiuniC2Z/gqATV0Sij/nSQuq5IwATJprt9vfZKIIXKzWTYNpiQ5ZgzIkQxCwmAJa+WY
z+8rG1a219F366M8yiB2VhqJSa4f3IbS15ULxl4b0InFOl+pSYYl5VOISmFyUeWvwlAJN/66OFPW
b3KKvQKqoltK3lG26+l3XsOZCmj/CO20xmhdJ5XBX9Ivn4ZbNbPKKaY1sAqk1X7YE/GOA41+5TwZ
IW4Nl5hCuCtMaGKfaQIwAnJ/ppJBdBijK/CZpxUcp8YzCtzCLK1ME0GyBtbGtEqmYUTkKZhNoPah
BVb12J3aadj5OtgxPKsaLPuLjZeex7ONE7nVP3FLXbLKCKt9CQNEptGT/qtlm/IbNppnTMikw6kf
55j18CYgFgY5pOZwYw4/ZNhOtxhdUdoi7A2bv7EE0NK4cC7Q21gdErzR0Tl0qp8Zw6Zix9C0Ohf9
2XlfqfjyNscnerq1bLCBIj8IOkXWkl02ncMoOaJYu5WlYJvyGK4HXMD3aInHa0hQxFhRlQ6ESfEt
nRFytGRnomKnCsHLlAa0g5rJ3PtYFDaeUPZh7DJQ8Vv/5nFLwZLSl59o926Hnxfi4mRSNjNZuttK
4QMW1MQejcy/uqY05V9aB3e4msWw+rIeZ44CZveA3b8/zAjcouiYc4yaFeYmIHbfiDBEvy1rmnxM
zQE2wGxi+PFpbtxj+nvAXIxARLm8xh9HoAY6NXKkJD/yomB5GU8PmWxSAv3DlX2q1wIK17wrxfze
3fxonCOoMCkxBvZVgXvACJ9oxo87S4VuuGQpIfwgZB7jTMWVUITyyuvpV5AdJNgBhTnsg9CbCTXM
g0Up3MNVxvu8oGKOJ+8ekb2iACp1uy9xEun7TEzX+oQOBF7juXcQDk3Relsp2iAIn8yP2CSnYOMj
qCUokGt21cZoqMtcavy+creV7MNsH1C8nPJ16lBYETACXhHivRIQ9piAv0tVLYviJLTeZvZ2z0ym
VDqe0uz1rcD3BxpaiN2uOnpL0XBz8XOloV9jqCQr/38F7+8Ysh2Nk7o2Oat2t8gIf30YiSE9YDO7
3hXUo1I6CWYkK/qMsB+UKw5BkLlcwO+IVnVb/RGQVfdf6SiTLQaszHQzUsb9RS7WT8m8t4kKLcXk
Aw9dhBmceUH6uOQ7qPQXlhS6Hq3XstikDTyF2tZIRFeHiiCgKOyJU9AvDfd1N5uDq7TsojxC4xZ/
ne7hrump4INb2sWFZY0hjPyEeeQNAGde6OdzVJrsJ5I6tpHz1Gcze0pNXu7XBVpvWdjCjEmUfbgu
9yITVTQ2rPXN1rXBoRzCgkxZBCc4wbx5rCNuDe6eTqRWp4WMxTmx1/Ma7jOM0GM6soXg3amnP7e+
bhtp9vxuaTK9oLKDiGnHl+sfXXhcxYVPIJOzaBvvSEhNlH7cm09KwB2rLlKGqKecN6M8F1ph351d
Bx87xhE/Q7zg0ThNRQU1pW2eAO3mXUbrpCjm1oHiIZ9n7h3WOH0IYTXooAVPuPIU4fAWiv0jOZnc
HaqQWKSqAS+87UOvSDLUC5vZ1r/9dEUQOUJI++0I2pJCJJfEh2O8ewIW7J4KMUC43DEw8eHiYUBI
EHeqe0hVGCYiqVoxscG6iBMzUZAjsfZ64ysDpGNdRfIuVl3apiVjT+urDicP2vDqhpTVhW8h2Sah
VNRKGaXZW86SpRmDgLBkAV8nbChz2EiZIgwhX2G7GfgykzceKtM3uyUakUnYOVc/8rx8544AQGe9
OO97SJQeFTgKbC2TuqPme1KiA5h+L28kJad/Jn4fko3AvGFyjccY9bb4Yj3QyntkGlHJzdwyOt4b
6a9WZhXCcpHy4BsFGIrhFQqJoVUg3fFYw1Qo9OM4FfMa2yK0bibTGv3grzMoMfqpLnV5XJYaWdrU
arLm2hXeC7BtbE4Y8PVfvC4DvnfcRkkA1SI/37g7Nv06oj6zILusfbV0s34rRbRLI4lH1ZqGY59p
yNCeAjCnRt3+PCRwCEdrTtq+Hf6VPpJMei2OFrFErhwjYzb979k39/BMR7gdd0mE1DP2C+6VCq9d
c6x3Cudwl7T9DW/BEWno6rcZxPO30tTpzcja66iQsaxDQjjNoE6BYSsg5vX6ZYpJB99Nh5zTXCfp
n4Uuw9x02r6W4nhn1aQ0E6QbRqR6vaWG/tgumnLa8mg1ago1fmNUhKqVO8N27nzM3Soihues0aTA
2pftaD+6+rqsMAQo83ubBZvRiiPZaUJunMxyvLQsR3Aoqyz2G/mOIGGildZT4iBPUJsM3oQGjZll
wv0zJC1e/u8tboe4D/gO+wEERuFJl+LVacS0UcBRFRRxmm1QWUSvJFfoVmB2Dgm9wDdCXzgW4IWr
WRIJXoBJof3nQ1reDv+NLZWuhc0vOyEWvJ03mgImFeQNH3zAmXHW7mBTNyrjGovy4e7GWvP2KAuS
fwnFgVXOG6ohpGj+mSUJWkSBsry+hswW68Wlf7Z99SRY2Psa8q5uwF4Ic+BuWIodEgYV3Q7QV2f2
/2Jc2tGi0KSj3CLq9tcYfp80day6VZe3BnvW65VrEnepM31BeR34lXZ5kU/8VZM8Y3P3qmCzKGfk
JE6X1+AZRBLNjkl/l+h1ndrBnN0ewfcO7EP6w3UtbGRoXejuxbKttENMMw/ayNVk4c/i8nccb48j
sBcHeKOSFjyGdUj2CmkrUeFiwQR6e+UGIwaBrwVAoO3t3UsT/nwWaaFy4ABbteWtQgAWf7pMpi7D
+BtAlEhI2epOs+UuVQMQKwTWar3xvb9pbdxTQ0jyyd3LBMS5jKHimgFmGqhoAskxpbwnK+LjlJxp
vLjjhRXaTtSphMZ8EBoQPoXe53C1Zq4j14zbjQ3k0rvVCaql5upmE0fXYjtLpHznJ2UJhanJFM+O
cXw02GRMOCmZf26sxGLLeiKJiqGlbsqsMjyYAq5aD18Jfs9uzDJIPQcN5Gb+QwS3klUcmAXSQFl2
ASdpddXm5VOYDe3tDjFtXYwCGKW0yMilhWDSJ3igAxTWfXX9FXMRaMORdsJr8UWs3xjlVp4odgJB
MDWk9FGZBcvFJ4JQ9pl12V3bEDKH5ATOw3mvNItJOBwcEtc5TYXwaQFu1PVdBqBc0q9WuVeZlEWy
yrE+IeyubL7015dvtkwuGa0GJyQMEm+a3VEcE8j49KM7lUuMIEFjyYSMNtBLmWj6dWM6OwFx3wjm
dc/5pIqefiNdOn+1c9reey0ein0HGCSl6CeXsxrnEFUPUK5JE9uwM0puxrZnTAY78SC27bZbTZr6
aWh7GY3hZNmSDlvjiEBAOaZMm2Db+r+osMZhBmyc8W4YlhvDvtECVb9wsa7WICfTKnsCoiSgrAjH
JXDGKkOQvuGIXcBXt3INOllRigGZKh7wjTIrvD9v0zJO7Hak2QERc2ZG0wlj34tQYV0lviZlLTEs
t9v4tzh8Qdv4gN9pSIzNVUNQMK8HSkRd9uDENRJMH4Db77Aa9D9aqgA0Fs91BQx1m3rUJoF4/E43
JcoIJXA5HG0a2YgoonDW8UVlkie7BoQ5zjeKk2kZiLQNaDQJKgiTXyaw0RKS/Q2L/z3+deryES1x
rdd65TiUGDOnnSwD1sJnlsREr5a5TUOk+OHNia9Hw5AokofTbjKSF+W38GtAiwSJEM2HDdqqQS3C
1iMOrthmz1h+sp7WnlXoa6dnoknFIIybTq+8Ki86OA8AJ4E6lG09ax5K5Bl6qGcr32BRayVTWYpP
wxopBqBRg7KZz0tHV9PKs+jjQHwsjYejMZGPDqu/wV7te5n81EXHyf4yp8cdv+qChP3RiWvwmfXH
tLvv7ZvLad0YX92PV81WrTmhket76dgGfGPl+UCuot0qUqX3AqvcTe1paGqgl8VndtrOu/GKwXbz
NO2IySVmL2nb6hDvW/Do/ATZWl0n8Fp4IseWugPeQmKlLdwk5AMCPLQB5lErKv59WnNEuuzOM5OP
FJXfpNTprL7Z6RjiuQKnGiGauEHGdzoyDTqB9XVyE26phDFoVSAnelTYswpU4ZjDDlkMyJfsVcJm
DDkatbHonfE2Nz/FNxsEej8hbZ6WtlvBQzHVeSdienZFPSooR/dUwcdgTzCr71Irf2o+nVmkpbYh
Nlj5aT2hBS0nHWAYfDQLLj9LFZEUR9sUZc9AU7M7tQ2UNUCPCMRraN3VDuWrPYwitMm/iJD0LnjS
lMF7SRnJJXbcJLhdZ+9iH3X76Z2p+MQ1AiXIxc0wgRYttUyuVemMNsJbVyA/6BqN5tROV97b2KxX
lo+7uMDKxmekRKbuphryRnyjQ2E/f6eh1HeUOczyG7py3H7ymFeWq+CBDXBxKNAYZfYZCs73pVMB
O5eHldrBZGAdGxlNL1cqGs/Q1sgelJ5z5j1azQoQ+yXOXbFxmSgpREuewKDQIroK03H8EH8leiKg
RF1QzF2m8m9oI2dTfYhbaHdW+3RmYkNzZ8XBgsBA4UV9WjEWL0a7pk8QOvDsN5GrbXqxZOE0P7A/
5365cLxySsrd8FLRDkBkKXijUGZ+xEvWMgtdFUhdvMIhRzzff04sqCTy6Yja7Ru7/Fkp1uWduZAx
5gu+l47FgG7koj4hnG9a8bc+OROKVCmg09zIlPdBFFSxQYvO00L1IQvV36P7eKausrJu/4p0en+U
jkzNjJNC7bNLX1hntt/OHIHa9o143Q0SijgZlRKTl893Yc0ozb7HCoSksBXeJvl4x+g57AKbRZq7
TVkiDwtwWpqZFdYuTSjLTJGY7RkSW/a9JHtfs7mPo6PuSDsXw6Eipm95rgHcJfG2ggv5OBHxChCW
O2Ri/6lnt6QwLtJFodTnz7tdPMnMg/6c3CBdKM/XDYhQIa8M5v7qDPmsHWTx/o3dH3GridEJfsdo
/4dX8aDl3fQfvSOb+17u1ymhtHQRdpv2yCXe1NJFjSKMkSNCUdEUYGTA5oIOQEYxWwKDQcaQ4r3y
U7jSEndJpV9C6jZLw+Ik8L4mQy/4igdSaSXdI8wnqcTUyk2wSA1PqJGjHR5Ox8fLikTuXylFe98l
ZabdSBH3GlWE7WGBvBTDFLdTw94aZaY3pxu1sRHhJcJCVqWTpE6a4FFFQOV/fAST/9fSdLbF1J6H
/sDDDzGe4/GC4uViIHFMI4FSOpVWB+ozHjIslAihWwq/CwpPBehO4fcYbxcuTaN9n6N9JymWRPnZ
sQQQl5k8a1h+NmcDPDMEg4k7SsJpjG4VxWdOoMeKStt9TmnDzR5zXyw6eVVmf/loT3muZB8Zsr81
aNyHujVvk5G9/F004YoKdMwZpb+d9eqbTxyO+tbA8LRNNpL0+2JkVOidXROkli4D+nhOpamCPYOu
s8tF5fSVHt3YrGU7HtR1nDhhXVKtOE5vv2gTxEaftcZAANSsbyDFfI4Tg1k6JgeWdm1775/7Zy7d
llmsP5RsddTmnRNC42G9T0OfSGQsZ6dQ1AtTgX1r/9EvbYG9IJO80peGvqEm8Mvx/692w0zsW+kj
ELtNfkQa6CsQeZnKU3F3KW2+ENyhjYeDxWSp1PVa4fC6sRYLxmZRtCsISKqEka1AwP5M8bmQY78C
l7dLnA8ZpyHvVAGA9s5LdeUNP2goB3Le3+f7Mpqg+4kEDhcS2hX/X6ApeaEIl0nUhewaWRD2VV5W
U4Rnxro1TxolHmIGl6RxQSHXtWaHs/mwUSrxK3V3AkxJdPMp6djn/gRUxjuWZaamFwKWnuglEis3
/KpLxgU/h5xwNnPESf2l8yCC8sw8bBQGySxEwKRho24ct80rn5xD2AqIDqLr08drNb1VM7DXOx8C
1AW23T7buXNOFZDAfSJZBcoO6QYr9yP35c3064Si16rwsiJRSdaN8ovFyTYtBw1RUAWNzypiBKAv
raNUMv5+FxvgAfq+Kj5fat62qIcLhTam7kKRBNxuX9OaAJ28Me7PWjl6dJgrGIjxyLDHlxm2GMlm
pZBdyyDx6NiQzP9+uLs2Soo0k1EPn4dow3PjPge8vbbN1bMNMTu0tP3VKbEcZ6B81vepHRkcXZIy
Q5ri96tLh5Keo2cyj7PdJfU21DB0NxatTTDJaj8fKKytDAaNoZg46DTddZDEwMfcv1kbdPp7pgY3
cg+1ISaDgbJt7SUS1afpiF4pugTT8nqj3ae9DcqWbl78l5QOIvPOAeM11hvEQM1M6QOQ1asCdf8S
N8YiTpY9//q6l4mEyb/FFzD8SayLVl/C0mXjORYRtRgnmySkIjw//89XwSZA9tVYRJhhinMscp3A
+5cWsArKqwOyMy/OOaWz919MR1IYZso8V7A8HKqEZvBat6W0O/2TSmIIg2xodZc+IdZ3pW6olt08
/KZHN5YFZCfFD5pn/WBc76IzFYTZw877ACAaWq9I6awOhV9nA7Dc4McmOD7o2eobhsz+/kOxVYHg
13eX1nML9uXyF/QMKKWE6TgWiFk4AEFaoLzZOdFSvvIthHBPflAHWAph3sbkYbNUc496nLeXcbfC
9fvYQdKpmHpIIviGRJcT0N2DLI4EkcAVnIwniYUkY+skdajN5up+tbi0Q1WNCqE5xR4CX3ZcbWbi
OOntuNAW/YHDnKLh9XwRiaMay7TFgcVH8GdUm94hMD9bottA38h26AaBAW8Xc7QQTVNJLzLvPoPW
AZxZSudnWUZEKw1Lb6tRg4JnhG2lXOzk/L0pMRbBEwZ9dO5yhVuwYKJvIanp9txcjNSU0RjlEQbX
w8a06slC7s4Lj9Myq+mNj/jQCK9v+oMhIIx+IuBm+hDekMXLVA7DyB2R4W3oSdpKQx7tQLH36Nxx
xWh85zwUwFmWAnfVtH/Vp/huH3WCi7dtvu6TlLv5UG3foyzxoMT2Fz4muqc2IUSGWnhZuZSeBCdX
w3uvRaxo0oypeFbbft0evpNrNO7baSTzc9JCH3iJL09EdHYlT4XTSrPBcagzqnMMPGl9fs9yDMyH
msm9VohmEUSMDHcbwauasiPi9uL1p8lsQW2yX+OIP64D4zaX9vAWOn9K6i7G4XlcjSkwt3/yFVWO
hOR004SZ/a7r8hofhSRaGtsPJJLQqRThPFsdV13wUE1e+jcZ1VBg8l1xYhORhi+Vi0aV2rAKcmT1
mHzyGk99tsHB8wnvzxbDJNxvUHAggrQhNzyfMmok+rHFxSBjQgW55RdElbNAx30+b/eG2KMq/e1A
OwlgYx44FzclHIo9kWbpRxx7iZuyj+NtUYTiEf/M56iT486qaIwQaP1rKglSmPPllLHs17wTRDUB
XV1WEyWpbBpiF49hHvlS7Jl4SVVM0mJcWHHMnm8WD+0aQCP2lnNh78rzKKQMpV/QH/oJHLwL7UcV
8eOCKWPE+g2gPmD55MxBWKP+f7djjssIwZM1zul3d/7H4/yPdkTmRF24k9Mca4mm72hZfjOjgr5f
ZgnXo+1zZdOTXQzlTN3uKiXZQ7FMlcPIj9qPYI1Oykz4qaF8qIdNX3QI2Hc/HqLnSFK2ybylJEZb
3kAJSeeq7CyxIedo1Zqn1XJhe/6oFq9T0qBl1SdLXVUNcE0imRSTyYNa+U40zS/R7NQBmmKs5TRa
En9kz7b9MBCIuKoxrhOk+CDe6uR+Ok9YZyk89iCrpKZFfX4ieD7zoXSoVm5wDbsvhVUSCpFuusLR
edQDsOWF3bAQe3cSjdrB75+WzfWy4SyWkRuPucHIFRwbVeSPYY7NVPswWf2Yc6J+IlkNuW2OF5gc
hezlEGau/UB4fCFEj+ucjEjo7VFIcflYRue/gbVYsbSKb/PSaeo87QTh7rE/eGxJKv6ELPcOmvKQ
1iXbU4Org8Dfgv+bGJkn3t3IfJE9OFIXn1NJq7rweQd293KhVGzC1XPzHHvFzbApYjUB+lPr13o0
ZMMVf8Ssz0k4Cg6Kk/TsmOLYRqQIKhTek+l0PaEmttPIeKUOfHnQcZN7Ifq09DH9YUn/FvBl93IM
ux7+89RbKIVwDKMf9I/ExsOf+m69yFOhAD64bIid6cwO2yvef2Vsa4qvYAq0CDN+bHzwXYKDo7ia
5rCQEY8UK8iBXy9pZ0UYyGRElA58RmLsYYjDE9JpmsmvcE1W3ahyxb+/6HQNMsqdLaplZjOvSxlu
gs7KLCfB5fZV9nJ6xrSuoQythjiOqEN196VHBc7SKXhnHRxD86UiH5/Q1RcM/ANv+bWHfU/TaFa2
41ujZ8hoP1wW5N+p9FlJYZ0fyUxxyESPZZk3QjESsQ+CeN0Cd2bSsNr3Ox6vLxsOcmHrd8LlaeWg
ku7W0fJD8bQJN4/nwSeDWQCAreFKq/PtBsdgq1aKOgSyugJa4BIWnUeO/h4uJEJKwmBjo/EurA9i
mX+2y+edr/Pplt0oo/mVa443he64pbOp5hYTg4/0z5Fb1YkrGT96NHb1qsEpO2ErE724gTvBb4/T
eB3xlZ5oxBUy0OeYqIaNCby8UmWKzCplsTybT0nWTz7G77R11T9GtQHfReuShvlzwSpHQiNDoKHT
+2VbfC8QE5tTNHoLAh93YuKVkvOpElUC3B2XLaTLKXMZtuas+c981Uxa8Uw4h9lErPmMKrScDomM
l4whBPXJfFWUJv3DSjlVxQlxpuhnRw/Cn+ZQJIpzBeQl28KSREVzo8zUYcxSS6v+gJayC6V5lX8Y
Dk947U0bVZlV1Gt3tXH/Z6H39iq+FJ4OlTrwx3hUIHsP6b746J+CnSTqC+4mzf0TRDibHAslSo6J
yDU7Lajgimw0SULIB03VAm8VgOxxyP2wGKTVObaDVoTjHR+WKgT5XI8cjPYeI3L8Rq5GVTbkxdxl
Dj1kXng4EBJa2Zi4QZPeQ9Khuw+XPUwzLwQ4lrc+P5NERwAgeyHtpbkrXoCYPn+9XrTHI8PxT6gm
bOT/Wr82hYgTIabTdvy56qvtEVyodIHkUbrWcVcdEvW16yVsP49MZOHae2U0h8Fv63Sz9P7Z0ntV
8Si+/uBk/LGyIB2OT4FURSADlhH6mvnCN/JbeoB1etYXdtLLR0rBhQlN1XbFWshxoLh8V1FHhP/u
uAp2LsllAQUnF3B9zSWaox1WyqC6Fhr78C1o6oZAf7aa3wxbL+OxV2irmKyFmGxgP/VSaZY2BRRP
Nc3WZgOi65hmNuPFYlgb2WXgCQBXmRsZZqSmIB4Ku2sMDMkDE7dGPdCByfDL2Q5GiUnI8zdRq3tx
CqbCaApc0rk18P0vHnJ8aohasNAmeYYzeWICJEWZr/EAFOauLYYXdDNNXM7Cky1Clov91s1p3Pgt
uZodO9wziIgKa1K3QTK4p0NeXtMQUSMbRg9TUF1Ib2Cf+JFEHwa8pKtnikzS2+9ILltnJSqIXA9q
tQg0JrFthi7IrEDAYJUcUfcrbVgiot8yhFY525UU/LXJXatclk8dx05UHm8KfIb996WiFritEuyF
DJzFUTbqV6qB5h3fw5jxTzRRFfqQ4zdoBmJD++RnbzcZmuKhbqE1JxoV7xWVUnSjK5AtRI1eSFor
L+Ij6dion6WjhZ48weF96mdjOIe1DENMPO3iZyoioYFNe7p2jQBu6DEsn5p17wUkSPOXSCefJkJI
TjMf1Jx2cdGJ6tJpf9Y8/LXgKwXM5raGTV09iRmYB2dNJsx6jkg5Oj2uaVxBDYCnoufkcXy9IO+A
T67k1j1y138xjSpdKFsFK4W7IWvPHpDfhSxOqsaJaUlIbKtbZrHLs7IkD2CJje2Az9/2e+4Ycsac
BSgb72/+VJRBc+iFJtGMshikyfaE9EBoKXSVzewhFM1prxdW3+M3xvq156dFU+qsTjBcHk1Tftxj
u1sLqCd1fBY2OEiqFr8kknz0Mr32D1bx5qwt+JeH5tTsGtGHAGAwJrgjGc/xf2JyrGh+DXFhsPup
WY8lVsTtkFJBMBin0y8viTxdWwUg01KWqnxLtg4lyaM1hkYeMDPKeeStKAVKO5Tv7BFwqmmwfR0f
Ro3ivdE/AiyJKnmiIFN+HF2sEd8NyKTm2t3bJlXkzJ8VCQy0B6skBtvIh8IilUBl8jv0fvvq8gsp
ErjcV96NoXKJE43jN+JpnLdAcp/GcsWun/GIOhowlvE/EkWSIV+DUojfGNGZ2u5V3RbxXzmtLwQA
+1RUBA08wrwaQXOAlUe1TeDS/vub3Zi3oT6mx2U8NgwunIE1X3WxlV4PQg05uTWpiDTSG1yV1R5V
sKrB0AXGcs3D97WosrxdJjcYKZGUeMMBgfaT6wwUSB5WCbwD0ZyXorjBDRgBa8t/hd4ygJjohMEO
CKJGwdkb9IjaHiT3jte2VBkyTXRe0nm5v3xJo0oxXETUwHpCBqzOPZDotE7Qa+wS61fxX3Ru5E9z
7/+fDAMwJZFH2FBSr2a5IM68K319LvYAEgvCf7L10lFQQ14F3w7KqJJLDEpn+lpmVQO4rqR9jgnK
qu7vc51vwo1T81Ls7G34hFvLac7x125z0waYKXbZvhPrlBuKq4TQcW9gr553XaUljIh51f07b5R4
vmFTPL137UAnkyhz0hNS1YLrQMXScq6i0QkLJGQIp8Ohq/ej+A6JO6uJ/+uNUj0mgE2SZZyXnQtk
OEUngAsWQ/xvbb2HL4FYOMee/nYdWdbHrGe00saBz9kbSpOhPoh6ZmvCZZ/75g0LDO211PZIKN0Z
c2/dWzEthIu1J68c5qXyij4qKUFPfWEU6NZ1bxpvUneaHME1UNUHQgqNk+UvqA1vSLWhzrOOMOcX
Foizx5Ov32O/I2rI4IoaRkYuAjdX6qYhdXmFmEcYrEn/as65Iqhez9V6UrYuUJisLRBLpDatrUmQ
4M+paoww4JFu0MnyadQUA3GHgJghc/YKBp2+vx/TwOEvXVTULLpcmEDF1g5aPw7BlpazRHHppdxr
jVsyfOu4wM6oG8Gv42WFvf5Ypy7ED/TPS+UqhJLZsLkaGZoVYAimea7Bfls2qyLguD1MQYRi1wMC
dqBL3Zos757PD7Ya6bz3cZdESb2zjeEoG9MN64iL8mh2wb7+gn+m3AzYOmuo9ugqaaKMo5if0ktn
1FPe3AfuIVkVLBxKIzinw6e/ebVzuPOCY7PCeEBd/Q8ka6iqc2egAePqISHHwExnVIWoBO+FFX4b
wHdoO1S5sxKumIBSGmjrkkwyisBCv9duZbLvEe1bAaNn0OAYPxM33Egp6oXcjk9JTCU2oGGXkS99
X1ljyyIkLzOmlQrI78tY0/dRJ5ZHi2xkjm8kMGOqH3xUoQfXwDe4w1LWFEj/qOqxZAF8kwh41cdi
vcjdNywdynYtdptDCpjLjVC4AHWl5F5ILInSOxYbFNQWLP8KX2n4LbhgMAs0/v4Guk2m9Dd+Lm5I
Xe39IumZoZeeSewiFHQMWY7xc355n1Hz9ib9VTxpO1F5Iot/EOtbR6mZLDgPEqkQcwtOQnoGXa8n
vxV5ElnCU9eFQbFjnlzAnITP9+4qVyvD7puAf7vpWPKaktGkabWgeCII8WV0kFDxwJm8UnBAd9sx
ZUAF74mtL2uQ8A0vb2CAeBLE7QZF6qJDxcNr0lJApMiuMnX4DG2d5dM6Nci8jKyerifKdUFCkcxh
X1FKdo4qvB9ih5csdMRHssbCTsn8fHxpXdEYP3Gpfco0/Te0nRuoyu1Ep8c8Y0ABw8Em5orx8dnl
mupHrnqMa7nztifd+Pbr576plckRx8hCVmO3kqfstmfUVFiwMpEtG/6GmYb6GlwNnqnnmZQqJOkN
94kPe5/QjNZvhiq6bjqY3A0+idA2Bsob/1yPIrrk7Xkwb36TyWK+56HCUozkji3sTs8YOy1RPlNt
tf2GLzaksjTunNwmOFCdFypf3GhpDPIWsvufi4RyzLhZRU0LB5f5NB+3FkoyzeyXtwsoXUqTP6Vj
n5PGDJxCsoVYjmfStHquA1NYdq9ui+FEMZVeJHoB3B3ZPCEdUXTFK8IEmkjG8KFyoZo3/eAWQDsa
YGiaRoslsFpb7xdzvoUSDmba/Y0a8m/Y3zv0rhz78WoqPNvDY+RBhejb8dVlXz7wy34KByjtlcz+
JA/k+dGrppHAW3wkUijAid0AXm53PcK57K4cEj1VlHBgBO1Qe58atag3KVB8LK8VFDCA3IZ9ziDW
q/QLXrRYPj4d6YzeV/OWTT6xdMV3Kub2QPkGhZOc/oQHT6Jg+tSpdExevMAaP0KW9bMj05l3ulA0
jnfG1DJZwFCt8mBCXp+MuvJsmWbjQ0503DWK9I3x0m3Gz0N0zDLeTCju92r1sGyCOWH/d15xunYY
snc1bQ40ZSFEqO2s0dzN667rwmlzo+X89GbqVoc4/nC1vt5I7oJ8FbSg/AOgR5eOUJaG9Fo9xkbS
K8IIk7wsDhz+F6keYE86+GSsP76I5NCfRUvqXRPkUufNBnc0juqEMITC2VJr0flGjZxIcMYwn0bl
rVl5SbWHEdhZmfamk2d2fWDNZO3wvwkPo/6Wb3/lP2L688SsVjIPkKKBhUYE03KDVGlOXvyTK9T5
3OvYCzxINAFihuEofyn19ipIWiVYqIAGZpI7+jd9DAPYVJZtv3X7J6ENpYKy8MPQTVu+aPSC9sQ3
MNJJpzGPPC3IjFZcxD39+3FixWvPWucOSZySdY+aH2u1IIkwN1It39cGCScPX+9Xk4d2KtktKEeM
o8akPNm8iYLiOKPbeaJpZ6RxQdkG6mf3hYWkVrCYRp4ZndNSSM8t5RDMY/58Lk/2bD3C3VADxcGD
U+bVy+1o3zR9aXnZv4mC13pvGpAFzTtYhld9ODjHOBlWUyqfTq4fZrcIPhtgjVjsIgbx54y/sRdQ
w6vUOotSwClwo4g3mHQnO9vcZlEQy0yq67nTjttynghBfHNOhQBBKssGik9oCDdSw8jKLW87dXjL
t3AgOXXKyuOO4rnzzH0ELFQ4wcJ/o3gKkyYTbvAUOU70cgtU8rh2vovnFUcbbuUOA69ZaZt64Wic
SGj0ZQ6YI/CvrLKmd4jS+c2jK1nOXGwU9NfMtlRhnIjDdI+UDKQA+QsZt5SBDVV70vqyON+MXxsI
lXa+M6Bwer26m8MqEOqEhbCVDXy/2PgpfuYs4hbkhbyCK4qXzgc3sjxQhtazdy/khLFb0h50ohGd
KVhKVgXyfb+BSsWbqWqkdVpKfGvypCj3RrI7A0BtqOrOTffXwVv9xpm2a4lcOv8YaYmOZE4qO5V4
w9AT21Ov1IFsii2jxYksHxNyHf+axD2szDnQufiDtb7GRRUx1+6royL6SchSIZopekg3UvXLJZGa
SsASJabCYpaap+cRwFLcBJxox66SWoYRwZuTec2XsUPgIg4qxC+7QQ/2jQzVnxZaADTtluy4BhxR
sttTPaPXe2RdK4yV72uJE1qZ++kLkYju0NL2U2uULbB38KUQBbNS3YTveeTMzgYdydMPk3gw1pHl
bIvG078ir5iZkQ/tuN7iCdMkmSAnoBLlwVwH3JH/vg4JuoagfFIbjokgVbP8cQOmnMjpdam6uDRS
ik37KVnxCfWYr/Vl9a83aMQiY1CUiVPrCAJxO91n4rUmlZDNzZ9m5ZZ89yyd4jsJB/wTAHad7Z6n
xGxRvkvr0LLoKNN/5PKHqqqJo6H9JzslUPHRjt2R1km5/6ixwQiUtOmcxPfilop0sc3gOc4HIhaH
j3d7tiD7ISm/u9gYPoI17U8P9h/G2HKM1SU0buvuXNy6iypgCO9KMS80fyxiBguen8dEnpAVFyRQ
OOyk8hywpZyuKzQDyzV6ZPMU+7W7V3oqFkRhSk7AGFRc882uywsQJ64JbO5iXPeXxJsAKAdU9xgP
r+ZTTb1prN2iIh+PbfuVgIjWcfpt2LFMhQakjRAMA4sv6CB/jrD75hFoJaXSkdXu7Rx9X/TAiepS
Zz2iHKu5MBRUzp7eAdZ4LwU3qVqBqdGYPaoRBTRyA5Ey+BWM8sx5V2TFgdoZNiCbVuG3/ITrtwJy
qJNgSHpoEB4H6/YUNB9wS2Wu6/8jQP85EqxiHakll62+Mr46ZEW4VlWHRDx6B3m2fw/QLn4pUycA
TL67hqdrQ3gw7rIUFRsTCI95aD9iNCTVKWUgDEZXKbKUiuw0WOZaxjEqY8XK55xzKLGklfXyYN1U
FGWd1L6YpTxfrVtl3d2U+kxMqcNbSMmRlYtuXq9oeaz+IY4u8Zd5NWe0Te0RgONfwkZ/Iw/QJD/d
QW93r8UgxxyAqXP8X36iST90Yzlna862vdEiYIOb8FEflym0Dz32ZM/zF7Y8VXuXRcQf2pz/njs1
OvNuFOnbMyr5el15aSgLIDFBDgV5NEhiBUGy2NjxZkorOA4sS1GSaisbwh0/4Z2r3wz52NIgQi6h
KI5AsGA3M/rjm5VrFaIhXRyYsAkScCoDfyH4pTIKkloBg0qQ9S+upypbQh0DWAzaiPuZzL74PRR0
fC1mxYbfyCYSi+mbR2RP5A1EskXfKUADaRTxtoNUmYp/B2DGJ8EymYu5korkavEid2f384nstt/5
ALwVgrreREbQXZBVcwrBpFUZ7Ha2zNKif7rnMhzXxCb3KvtcKdDh7llZvYDD53qjIFH00qwIb4fV
L66oeh53hNo1iUKah8fhXyU3+F/Tv39LpBVPiLkDRmPvxm+As/fa14zs5A65yvDXqjIumG/3hTVC
ZwTAlqN3JZ2sWIiMNmQ5ICe97aK9axv9ie9xUSLuI/UrCr9byuWuN1rXIn8mft/wm6NgTH2xhj8X
nDoltKJj8JIz+nt4PQgP2DLYqivxRUdywgrSYUUYGiB0f/butYel6CcDgdhvT7a4WHG7SLy5Taeb
RzouM4RZ7hUWp1pgXn1n8ounNpc5pty1xirtN+dgxrvKw9LpNef9oitG481OpBvcx2TEO13Um0Kr
T8bjFLsn/nExuxIsPxucdCQhmCF983gRVP42R5CXyxwnLFk7eeWTopXLiPboGwlvLzkvglvxiP4W
xiT+aEBKwDfDvToTv9O8qZtL+M9npCztyY36Ns9U75ZonPr3lJdxuj/C7WK6N4VTyzl94mnFJ5Fp
ug2I9wT21fUhuZpQzzZWI9zcW3MwIuNVCZPau0FmsuAGUoraCf/PLlpniiRO4zoO7ideOuhG/cU1
tSM95Re1pQHx5WBwH19HllNAIu9495QRx4BrnjGJn8LVzLALa0Yk1tR/aO5RkV7soe6AMorx5p4J
rIXQ8wv5TlNArpX1s2v7wUXuXDg/7VJDtJYIIdg5I2c8UHHJJCFL6NJENxwnwxjltS4zFq06Jba+
BnlLe3Qj0OBeBlmI+kA0hfRaJ8rwHVfvOmbLal/TXA4dBhtYg1U/VatWOfE91GdphovZni8cJ7vg
aideXNq3ppJ1DrQIteo21Iual5793Zab6L6q5SN4qYTIMUWYmbL5jDqmQkrcV80eaZbgEEXfGdGR
S9fMecvB/tLfp90ZkHiSqMnpC2kC8ej+CwE21a8ay7B43JMFED70b+z4lUapFA671MIqmfys7AG5
i2dJwOqRMgjzc+93QASkJx/A4cCJvUKuQV0BsZuhgVzgPcbC7G3JM9TDI5PekKiE8101Af5iAWpz
xX27Jd5jNz9djSVwydYn9meuGHZVZZICk94LVvUxs5XHnfc/q7BXgADHSpvrv0yQjK+zU5HYvpW8
XZasgp53onHAlL46+5VDFmitBrcif0h+ajKN2gS3aex674UtBO9V9WKJnA6gdCobPQg/fA0b/DTZ
XQ65S4wpExNzk+YOgb59+V/bTJTPhFDbM7T0Ul6B/RBgh5zcPCNBmplJw0PtjOGGhoQ1BjvAR1e7
+sjhHPhqxt0hEuYN/uKseYjTSdnM1PC4v5W1xRG6pnYV9dwE0Twl8dDXyVOuXLSULTVFAmXw1h4T
pNcETkoY2MtiG5fLgc6tF9d5YhOux9Juro/5quDJxokQNgGJkFAQuaf3xqRNbUHL3SgrH+2pDfv9
uQ2AZ2ibAAH28dD1gygh1xis6wKmBQwoUtuord9NgwS/LbNRYOJbVWCCYwpwBe/YHYxynLekYvmx
6vMVhSyx4OEh/03LrxFYDWTGZx1pX8h93EuswObvJKTFrNq946qPK56dphojzBg33AnWxQCBIOaS
qE+HYBXBkj2vZG6CnQt7W/v0l1DLVeIz9lLoAoW3dgj4tOX6V8ZlGZaHSQj1hZlpQcG4mGSmRWO1
K71JuE9sUNZIRTYHSVZjjXLRalMoVarmBjKwgc2SRYqa28Bfgz0gYOQLFgYMman5Prl2zZLc/guK
4lLokULfju23NZH0PyiG8VxiPmp3PamO5nbg2p5TOO6FwpTdl8m14zByaUadrs63+hoWaYl2NLLe
GNO2l8m/qZigdH+BlGsStYJJkQ75c92NloRFLPYEAKdCJ8K+1aXA18gldmTJf+6kjm7kotHhLBUu
onMjC+ru7RcMtMnXWrpu/OeA3ASVhUElDcn1SEad/1SNKhqb5CCLmNlCldybiDcQZSDXmPDE13QW
tQH+UeyHDtRgTTdx7rRdRu59OlRXhHsdZM/GYn8xCjpMVn3ooLZbXiRSBkdD90ZAPnZ7amDOs4Vx
uc96egen3mEArDE8zZH5c+LoIb3VRu+3FWJzme+BFFR1AdxLHiq+P7xB81/fiZIY3xmy4fABfXJJ
buVnrRNkMNePNgKfcPmMEbXOgzY9PQzZ2btfEOT+N7It4DMABRczHblHjPy01K42ele6R6AByjXo
agHUgEbftilQRf3R7to1lZ49OQvBdZgziNo6V3X63Jasj2ZJ8usIKiQ7hCIJ6MIHDrLqm/+Jl9YV
1FKGKkqUroYxdvHZCz51Wsk/8OO0Xtbldx0e3eCu2yQy6aRC1C0ZhwyQV8JE8jiOnqTV7oqaagIW
wRhOjLVfAU/jJh63pfhIuz6C+5ZD+6/rJKcCudpikOPRlVRRQTx2q9LAsq1FV3OhK+AqJQyd3GFX
YmeRr+dWhGE5ziXYoLyme8gnD5W5n30wgFxbvM+VoQQxkrpPq3Esnr1QHPfOeeB+vtMmg+OfWhYz
/pqqkoG46xJAw4gEK3CWVYlOtPgqWkReM6RCLbqgdnvNWspJlKnwUO6sKDHkI1wvwv4YeD8n6wgB
zhmnmp+0o1BBpe2VbpB5ftk/TjcouELWpTQhWMlL86RAIotdR0yGCKxYaGhPsqpZp/ZSR6I72NzI
f0jopXU9BTDwmTgxQb2hc9hABqZJCDfbyfNrGnlfiCVdFj71M3i5sNnXQrQUW9M6wfa1CqGN057E
wejSW50avmi5N6znWSyqOX0vIFWsLRlhhMw7THPqyMUrOJQqX7s4SLGqtts6i97UkDcvDk6OTXXK
4KdEjMmUOCjxLSL6aiauBT7sihGTWla3B915+N8IP+4LY1hKfh7MqoxAg0mZZUwne7/XKDOC4Wlk
Mu8oiieOUqcXbSDvJJHr7qdBEPbwCy+D+bXJNVG5vYp+TI6peyYZoUspr7vIo08PedNHyZgGk7Fu
qkDOxaop+Rp/85fXRMWlTany8naOcmTOj9LcH5QHSKrThlwyydoIsbBUzvPE7YTAbnFLjIiIpLWd
bCFdu29sLbiqG9dupJSek70G3VCbff6m9kPr4Eu1utOFL2fhRldZoho58n3433UuuIxJkbCRiCSF
6CA6W0vZCcj3YaiBDOlfkk1QAAHwpphfGxaHYugaDitgaV3lZiZoZgcgJgoAJMLgDLYZu9Ckhc1B
f+cA55Tq5AjAW4Zq7QaIUZPwFtQZs9IPCndpbNucA177EjYswwJmqwHp/QioWz45kutYoyuaAkhg
W1S2selacDohV90Rkof4t8vBcRtsJ9IL7xKCPgl4TNtTsBjLN3WvnvA5VfPxPBOiEQEL+6iL8+se
wApHy82gS0qovBlmizNXQttLKgWOjkIK9iSMLKzBdVYhEE+ToGrnNCG8aDn0TtmP1nxkXSUDEPtN
U8x9Eq0hV2/nS565i1YjI66Cy/tM0HARZUSdlx7y/zlWxn3j0zqs0DHD2X4XmT6Grgtnmtt/azID
btj2I9UdQw/5PQjQMaEAx3ZQE0yACr2Zoeo9LamZpiBGiWkylJ3g6C50oYQxGCNT817GBkuDja5J
5HBLI059CFnuXFxiuHKRG7+8AiYdh8yZr6dfniggb7NXKY2jYt0H5iVRb+fkO5VzTQ6rA4o6A1Bl
DeWr6EbL+KuLNqCXXxbTiShe7dz8E2Gbq3RwLT8uBFsB/vI1ueZUoKNs2cOzpKvycJvOCDmVfUMz
ZZ4u/+lK4BGBoXky0/6B2WrsiNqSrOIKLg7h+5vssxl9MbTXp7+BxK6nSPCETl7RPoali84HCIii
+YJhEh7M4Qjw3B5DPe8//NTOGT8uRJM0qoROd2YKfIMlBe6ienBPtdqC6GAeiG996jSj1bumoecn
4e0/mXAgyEbFx/r0ELTcqASuieqw8gPCLGGBg6LQbtVcaBOC7MxyGF2BaFCM3c6KEAHs0GNdxyDy
oSVTg5kfxy/NZzFT8ESRaBSGocWLoKQTiHb1OEEHLrLEYrJZd+BdMS2N3djGt9RN0pW9Ac2PFksk
lxydSZwUFAB2+b6T49T/zXUT4l6vrLkv4lMnLTIeYmKiyFxJaucjfSkpjMy2dYrsqeka/kIr5oVI
uHF+V86LTQOw6G8usuLiOY3lO/lEfA3QxRGzxjbGMJhty7bEzIk9JRGZIQlGdyqqSVZtisXaTuLd
8R/vT/PrlOtXktRhgTMMuxuzp25W1QtuW79SqCzLXQQkNadIbnTS7DJ5EwW+qDoodHhh62lnJIWW
MloAd6BoRELT2JVIZ9v0Tp8pdILQgrxgDe9/L1WECVdt9UkEgr1osLJ0sw7wtAiaiPj+1sq3vgnw
G1i6bTNXRxh8ujdR3zaSk60bMwqD1ycQPKOB4AHdskMrBqkod4UTxl58/xWDhKSJzwB11k8nLwKE
yv42j30JrOpPgTfnyVGCf0DyCZbcF/Rtpjx2bq0dzbFdhuICs+DYtksWCognlnLTfi+xGT8hf6aE
Ddrk2XWMh8V0a/NEtzB6JW783UQC+5hAB6sNgovp45Nqo/pDowmrNJ4TrC6J7H+Ohaaom75kEKCL
L8VxfP3/V7G2DxtGYxygbxvb/GrjFkxUEB9/flVxByVWW8lHfVGsh/o8W6eUJw5SVJG/GHJdJ/eU
OwPM8VvY455YqMfeOa4hCREoLSAj5U1tYa1pfEGlwwXfG2NfhKYdmxUHIum4UPtw0YulrqjoeKWd
S21I0yPN0gDVHXp2DI463Bkb8xjafMltES/w2zYa9BVWWU9CNoIOFjB9ZIaNoGFNbz8Sa7o2qDV5
3ZT/fEmhc5/qvGeYn3vEcWKiowKuWVqkxQeQ6nmRDfXvv3ppaxO/YaCkSFSIydu+SO8jyf6iGj2o
kz8NHCiqdVUmOAmhXlfOGheV4oXRKnqbCU5Gxm5tlxvLk6VrnJcFgcdVnOLcKzsJXsdE/Cqv5bma
Nx4keYvAQAsCKvH0wsw5nJp8pHZK6OjjyHZMbcVU3/pDYf5CQ/jWwgAWbuozawsYz70aPWpq68Q1
ZRLmeziMDt181eI+VziuquRt6PLoQVo8z322EpLMLntuAzHL/LHO02En2EnopWk5wxtRyWYPyLfa
FjvWUSgh0BfGO/A1UJurAhKy72COUyb+sriOa2jFHzIvROqeqpWoVlBGX26y0ciPUi1i0Scv/si4
pldytrfpTyEOQHUXCLUO/kotDiOqYUi9SbzKGNcfhTqM9VMynA25dzsfBiKFAI652WDEMeMQVhE4
IDJH5siZ1UC4cwcymbG8uAoLe89dtmXk10FyYg4acVs/Tl/wfEOAwL9L1kk4sfXDdsNaPMDP5Zbt
5TgKKTtmGnHqHp8ZhZBEUtR9mEsDvCoMUYqLgmk0NGhWOWcp0xCMIfYJ8m9lAFjXLPqmFnPlu6t8
1cpjy+GOnRJcQ9KsnA+W3avRdOXjJDNElkYw5sfS2LLJmZu/hSRMTQU7dCAIUlcN4a/k7E382L45
ERfvveZ1FhKkxLF4HkQvL/k/RJwN7/Xo5eIEkoWHaNbKKq75HfkdMcgI64VYQqktOLcrIpP6jr7I
g99YAF3kDM3S+1wYsCNykgBD0hzE71oA7vEcGCzcbvyeCFM91Ge8ngEPxSuzbWpLDywqzAOWkTBE
BvskrLkq0ZPsqYEYOsUgL1qiBE9BmfKdQs+0E02CXKs/no1Mv4iRHad1MVBA1Z5RuyhB26Tn8OYw
HU4WK7SpFQ+0ygww4sxex/sqlIN5FVlP+rM9T2bwNIj+Y2fZzW7zvM9yC4dfkx56r2/uj/xMOIQk
MZZTTN5Ck8HdaXr0UZYsO3VHWhzerdAy1+M+uWeXt5pjMOVoJDyjlUNB4K+K9a9fGx1B/PRiu44n
bAjyJ0yiGIb57msCjbawmKQUoOJqQPQ8ELLBNhhJt3Re5fgHfRM2BW91XWjMQ/7yci0o89YbUTlV
5cIHtvNf61rrrZxkujetsUi1JAz3os7MtU1MNVcm6Gm3XZjLksMFmc5aDTOkSMjy80wSIZh2Zhq/
Nosfp7pyswEj84Ms7NgLIL8cPyw40BrCt/xcbQBPPFM8KBPPJCYwGBGeEJ+VKNRidKy8REY4/M8s
5p8hAQM0oBZO9+SsxZC8teskMMibhmB/8hti5af1T1Gv81v7QKGFPLsBHbeUQyVVXSkvZawZnkpX
HnLep6ENVGtg7Ib83lxUD//E8HMKAtd4oU7WIFUdjr5/tzKVre0VRXR7+7K12rJCWZFW43TsTfkt
qElJAkMF+Lwjw4N7Yk2latThQ8ByQiE7fhdJlveYs1UoPUZClpvycdIKK5etOPg1eA1oprhR6Dn3
JgMax4iwyRGEKV81fTW81TwzATmFVsYRl0pP5nbYBx5QPDxY9N+96HXRdpE/6EYfzZ34ZxJGi2qs
93X9y83UgiULVUkyTFjwcR2vfqMSeWD51+TnkLtcj+6vKiuucDz68CyUpqD7Qr4j6FB346SNdS1q
nl/JQ/51apfGjGcVnlCrjzvZRGzHTN/n+KFnIiHjWvtonT80vegR5cx/e//pH4HbAfYdixNWtKOY
AdrcK7sqVg+o6ywbz6tUvBEOEq2CIoBdXhymQ4Z5DxbqaTsNO+Tip1oOEgJ+unXlIPEUW/8rPhk1
96bAxPDse2QCL3UrFYDto2MEMeCUgYZ8hWAoMvkkmdx47q6OqzDBIbEZDXccLRckTWdqyITub87i
VGFkoscL2kjWqah0RajwePX9jqqExiu7Q9tT4bljq2vVj0JDcuDM2L74hC0EfRBEnILDpiJoG7Sj
pmTY/AN6cglM6GKI+mpQ03PAlphwetCLD15erRTah8xxJ2YCXZ75O48tXzxcc6dwWpGVYwI2pXC2
T/btPoOOOf5vnB9DpzvI55h2P4VuBWB3xDXh4QJFzHX/M5zjI2QV20oG589cqATgdghouvsRWs66
mcRrrinBnxTCne9ZeBeHIDlZifiLfXhV/fZAwvUnH5GPOfT6tNuCJxAWy6CDT9Fkan1e/8MZJmry
ceNuSLR48fLA1RPNCyZqRwIE01rYP5gTehUQHKat/SZKaX/AxXpiKa+mHOzrpaKsAeO0x+Y4FqLH
zXp2xX5d+MIDQbiC4ojQAo/Tp5qF2FiaxuyN8KjOrRVW4S8OxUpMrG3LicV3/+2f68iij0BQFRxf
bt1pvutN97emuub4uZ3QQFLprC0Yehi6NUGVRos071FP0G/b0mzvEUr+vb1aPP3eEyRYytepFAKx
dS0eJpdrBZPquQWHt2Ile45cfhPjibTZ4Ratsi2ymSldpj78SAkuF0nyDQjiuDh+OtSFiLsEXBWm
/Bs2w9INWYpyNu0I7Hkh3AeADxwlf8sX7BvytGFo1SfVJP+Vmh47SN5qKE1gNHUWDi95X4rTt3ty
i8V2LwFqd9ewSbx06HubdY+6dWxsqgSBOEKDfOHL9O++Gkdd5u6Ba91MxxTsRmgj6nogy17845Jq
qNHHNJH3HV4DY3szWtuIMrM8fd5pmTFPCGKrpoIAYyALH2GM9N39OwrWbu7LSdjqzZWPSpU57CVq
TTjxe3AQfTIgDxttD+b2jP8h0TgmnRCF4y3HPyqSgmloeYiujl3Llu2DpewkzlxSeqswNAE/7wav
66jeBLILcETLBMD3pbFX5vU4SJ2FlM264x6HP13WPudHbj4aRaFlg8Yjq9CHBFmHVpLVg6QB7zOv
jVAsZo0rgcdgeyPYzYoYTNkgITHUKLnoPSIzK28wughIr/bgKabtzg8PXAdQUa42i86Mkqu0cNNA
PkNruHzuuTaru8AkFPmz8RKOaBsh9lTti8kMEqyd+Y5kvjhurRyhOQ1J+vo8Ea6FvDtmnBXgzpqk
PsHTcya8zXnVfIejZkRyHKIswvISdYFkRLQ0DanfWEagTa7F+Ff8lb7sy6OvsrsXkhYQT1pEkMDL
jdSpWhTdec39rWpONT/w2JwOXvKLXCJoZ4zykmXp7Qktpw4wzJI9VXIPmH7bYfEISyRwIRAW8M3H
U8gMlcHnekMSzIj0z+0+HwZwwWYNOAKwka7G6NV4A9lTJa1IVap/Fy9JxmrqptWDS8z1s7vORvg3
fqmzNsLmCrxIYkeUo6giA32KpWXxjZcl+tN8Uy7A4lVkM5VD8b26CERz967xpYbtHGBY4iDmSZSU
/Ezxug8obPuwOK4OynyVsbQTC83nxt+z+/9Nb8kBMKiV9R9sM9z0cbmUdOeF7j+4zlpoyYaBHOc/
4Qtrs0cUGNhww7ehqXaWKc6K9hrwdDkjhdRf3zgXJkd+6B31VSHWC76w7Trkrfo4CaNWDRnoKHpc
6Fj0AP16ABBE5fWekaZceerCAo4+/0V8VEw/HIH1Aq2zyFIRXnoYf+G35EoyFcFshWRzZYYvioL5
soYixV3sR8mQkzlLfkRHaJ7gIWLMt0hNUh3bgSpSwZu3pmLjHW85Peugj7oCxvVznc2GMta5epO3
XtqCVGUo7Av88LRtswQffxyoNGzuRG2uCBzqwZ4z8iuvx7e7LkOBMyj6mQO58XGXg58dREDs0NQe
HnhE7Jn58pyOl+nnwGsEFABZhLEiEjPu8emnctAYdHMKzqPycMBgQw481j/6+J+Y09E8y3pFG18b
LlP5RSJ0zFWyQgJo4RbfKMyJmY1eMmNsWKyV/0qHCx0/0R+rpWHI/UrISHUFTtDdVsbpe1Qt6DI7
mNlSKsK5jjU+FnNAUq4owdJsofGtKJfkNsrS0j/nM+x1/30rgEbsUGMqjll0hjIny5/TZLBFlNC3
VYg04Rl1ZOx4SJiE4cHdSInwggCG9jW/Ta68yc0K8MIbBhrS+nuCA/RiZTvyHGl/URtjgmwTHeXJ
hGKetgS+DRE9xPdJBrmhj0INsH/Vym0q1d1FycXqpyfS0UAcbmBZbh+8Qpw8EY0RkFyRhtOonrh/
3VPPgUyH33qMhcmdPbBm/g9j0w+0H6FrkYWPSgkPcBpPkL0NN6yCd6XNWLuCIiH4FrwqeGt8Ucw9
J0ikniy8u3vWnXThkCpfLsiQQ79639jp1UZjWV0e2JD6QLmixpC13jdPmqV4vPt1QN79z+qvJeTT
cTvfE9pThKdyNtdyWS8Yb+13yKKEFVlfa4ks0P/7w5VaD8cFnp1r+fJgPtYnWenjTMKLb8QMNLFh
P6EjBihheeQ2MnbtYQL6nB7Y4SvpM3GzdwuwqVy2SbDHDH/LEFb96ALPZ93/jTtwEkEEe6tg3hHo
G6CZCYHoGOSPRjvOXd8/sxHvpKO34C7/Mfm3yF4+zoNet7/YVOZCR0CYuRwZEjFedCLX0uc1a4MX
dtyBXoQbKYcQVxWqZdDut84zCi0EQTTmW3FeSkHkJMI9QSiEbCHtGsH+hqG7eJlaFHmYqXtgPeoY
OFCXeYxSysIjr2UwAPU3tPKn3Rpl7nUlGmDqilFkodhh1a/fkH6Cxdyq2MKz+7y9TTCrb1SX6rvF
exBF6d9uS4DoVHGNuiSs1csLRksi8tKH+5e61FCb3BXfEkcfYoT5174tjMBSsSun6CjBjFDCUiHa
rQ9pJk8n98dTttC82ByJ0O+YHDM/+Z11G5NZvWmfBajZfSj+g+FduxepVSr2fhyn1XxNAX+dF+4r
NjZkNq50xr1uq4T1ZChiOlCfGRi+H7a0sqnDZUr976KcpheFlzfmKbDINey4L2mio44Mx7tkKRek
XmnW9cJAgiBDPYPXkfZx8yE3vqobYO99oEkCvQwmAeAwNZsyUb392K/K7jqFTKg0WIb3jDIcS9Ad
1tPQPCX+vq5MNLqivSxi1Uh/GRzYcsaNyuGdgP+uZQi97p42Lscn+4iO0eEiUUsWi8ZAN5Pt0H++
j7sztgFaRFoUNHisRGf4VpCsFla/f/2yWLXLZPYlPIVguL6QEU14hrknD5LaR4VHFKATK6X1rKGc
ZpNX2JILOqEjL5+eajcx9Axpc5iyaoL7//nD7UjidqIhiEm999xxq7WosHCM29t2unxWUb55FsRf
LFNNFsJwmKEIRPV2Bg35PFIwSBSk3+gM7QkfFI6eEyAXLgmSnHjT77Y6yvlNTOLle/SKxXpya5r1
dRHVKa1EuK9G8/5quy/SLU2Bye6fvzJNRlzrZW+8+U6QmjWvVxxVGP7s5jKxtTn5b5e3nf9ydpRm
4WfJ2dMnFEZ7Kd+h4HZdnqzp3/IPXLYGlf51A+lqs4KrRpgXMdv9Vm7I/p4yMIPGJv6HJxq0Lfms
VUCVSx9FqH9HyAZ4PwJ9wOvXY5OLlqNliy1l4TSe6bdFRrBxNwYeM3R/f0GiK8/TgAN9Y1aa3Wl4
TW+whMgXXGxkNPKlruxvU/WGq6RPjwuXKa3lKEYPceNEwu5SXng+GhS1AJiAKd7bYKrh2MkrAiOQ
BakRPUemmhJF7vyzp61eHW3xi0HL221/mcc3dQAb9oeE3slo8upIRJ9mfPoo1VaDqkrMAFPxf/ms
CEzaOnQ56f2LQ/eA8Ti3o4skvKQcUAT1pCk+lthtThs7yP1HGDVh/Vus+UUVs7GCxS6lPREiIiuQ
vB3mTGl663SEAH/u/N5vwlvyF6lyIrI23bMOwnDeOCmjwRKCZ3hqZJcWr/bt+6QSScuSNPLo93IB
Nn+YVCwbqZPBCihJsvIwupYzvpS+vYuhFxOW9j1nga9+TiFzp036tdaDl02jx3u+o1Jp6VgikHNg
fOHTo12GjnZipQ4c8+MhlypKOmBFM2rEpqVTyQY/rwpsIndydg/GoQGs/8oZEk1StglvCHor/jrr
G+8Vtl4s+ayn2ReNPWUA5QZjuzv1jjE8j6Y1c0WcSrlSg/GUa2ki2vGkQTig9fCyoy4U2WY+Aa/J
4iFpRlIdtkb16O5AOe0OfnC6Tlo3wlSZnq3z308tbUtW9PQIe793tDeX9RSThi4LUxw1J/iwsyaX
DcCYxOI9UnC4M5vj77XabP/LdBZ5rcqF1CuZ+PDUqqD2d/KGqNqMLy3Ak4oE75SJkuXlzR2Q/L9t
pfWP4c1qfVN0np76M3hepfzpjlse9AY4lsgCkYtiKVVvjTXibHxAQXtRfRXIgrkXKARlvqQJXL9l
ovOILh9mZnoz+h7z6Gp+0zjYuYysf9UfB8bctuFG9lE7SiPpY0hCQKIxMwcHKZ2IQENvKTlxSXQk
PGfgop4pLksxmlGQYZa8GPwTPcMrjOPuzjYiKwRPtDUxnkRsZjPFpN9GZB5OK8Ut6yhFjeg7d5tY
QHV5iTlhboPff6RyUMVljUZl5ai/Fz4YhknGNjFrfKe/zNVVw90nFNFVP1OjSpNodx4/BzskpmDn
9B4+d69ChrmBkEj/INI78T9yTopaxkoKggqRCL20VmldhlV7ddVI6r9Z2BgtGp2hOsvaC4hGalP/
/3nowm7xh4COrFiJzDNt/BU6EP54QBO3gij8LtFrvSyHsav5PSVfZ0JLBjC/E0GTyQILjGwdrn1l
n2wtHMcw/Opww4Jv68BcKR3qJ+z6dGOQ93GS3OtW7nWMWzIbTGHA/wYf2+HHlFfq4fpO00JiMDjc
PwBx4NKvj7Tnt6CRYSR/cu3z64QBjYVkavsb6GWY76pjxQFeKp4ehTrnGM0fIQUlSzYkCmzWx2OQ
Lz/IlJZU9Vmy5Ec1vcN3TVx6L5tOfXLpPYtpYCe7+oogAn5MvDGfmNozSEGVY2QWLtRkusV2u5WJ
JMqXV3dcaiiU6a4yCHRXoKq2G8wkoPygxc/coTeP4SIFLSwFY3iqmRFlxxmIMmsCVzhVbDD82uAf
lA3WOwy009hOhIPjSCaig8gfKH8u/gGrWguplhd+8V59Q8/lctp+lJVGOZdiINd8mV9xMafvndGF
mWlnDkS9BniOMGe8qYfEaHqZPmjec84nyCk51W5GSUAz4drZXXB4kZ5K1IiZW4ArdAYIRzQGgTTS
mq2N3hIU2mgXFSrH2+cN6g408yeLlKzTfPuX09v49tft+gVbKVUlCaPGFknzyOWmhue3Eo59UtyL
BJa5jdhBVZkOXAx/tln6VAolEnhQrYVNsrR9E5bTw6DsuIhIFh/FCH5ecbT/5QBxyOPUMPpTHQrM
ftKlfnx1ogu/B4RrC+EzyroQOqJOy+onK4h5FqlrCe6AxEy91uXSGp+kXUvXPuFiQ4QFcBDfEsRy
IuZRpxO91RlH1nJNHv313dtu+IhKq9u/BY8Lzi0G5n8z/+qUDRD2TFyg9P3bC1Msqd/wiKW3lnZq
K25o+7H/fJf+aFq1t3au3e3DUkL70YzPdHNI8kIGW+g81amCWOaLybURnIb6ImDVnxMODHXuKGwD
brtDI5xfpdKEVv1oYxxXDo0Kj8+Yw+Zr5t8R9RyQ1KefDblmriQiCLl5RhtRCXmivnuX+3GADrAx
0oRq91lxWltdKFzjfmaS0XKjtHSlVS1nxJMtswLdJb6QyfxsInQWmzokblL72jH9Zc07IERiyipf
I3NPHPtr5ksY9HzFytRAAZpaD98Q8rjlkYb/eKFbQ+GRngeZvgRNDOexWVcYLKpUI9FjAqiVjBdj
rLkxsEquhhV3Lu+lq2JjWjsb8Lg/kFMMM+am49sYgRxzPVlv1CH6PTc4tRVrgyxQiYbobOGseSNr
liHCQBPuIlfKyhrcSTubI2OMMsaL41X3CR9+gIjxwFkQTV/p6rEagXYvRE9u9USO66vf5bKNyHG8
Hpd4e37r9CeT0trPtqBqyRvllLzCr2wjq/ROZY7n0U5cmW63lQaQ9XUOV4/NJZzFzglOPiR1ysHq
rkMqFljPPb7YV06yDEuGzDe4amKBt66dL78Pb7KbcstOdqkIAEAReX9G+Jt9DrKQ4zpZ5ZjhwAQo
LBaea6a/UTbNURzjCgAKmvcQNzGzoijrIUi6Rb4XNrbY/G2FNcl/fG1wgBrDuhR2vXNF07ocFIPD
kKmm3js/NwCEUdFuNQiC3KLfPXGjaPj09sCX+oogCZdXDXW7VdshQSyTfQNmYCxWJGR02P2jLubZ
4wmspj6zwEytp0giqmEIR/m09/QNNMSLq1Jj3mW3ln8f8jXDkDmKa4F29b8Mxdt5GrEmGRTIvVt3
ks6hosE9vJ9peFOdhZYkSX9ujDaZOEb/5diAxaF5aFHkqSd12/OHLILyiLCe5d8o5qT3WGn7VjQp
mNf9WbA60kA+zRhEjPTSGfNEsEBxamcaIxzVbQgfjhXDyE9BvCRRtC86hwG5czTqGX7TUug7fNxb
yCHlIv8xFaISOle1HwUfniR8hvrlE58+dcj5Tj6B/82EhEozmXTpWLTm0LX8IWbOcM3LNdgfHZcQ
0sY46rhx8wDIjgxSBKKzuBb6NLyJ2wq86O1B5mp2y1bC7hAfTuoNlkdnftCqguKyf7YIGIaagzVq
JTfEqQQ1TCFByYYJLiKDrJQPvq74hhOcVyptxKbCWQGerSwaL5KddNEXFTld17D88KyvaXpBSnV3
fYf8kEz6e0WvxMtO8Ra53Ah7944KAM0uUGhhbNdFtJHZT805qtdelEslTIvhek3J/FkhzQGuJBSm
uunm5PbB+C+nBDrxGfaDiH6Mx/BdEEQnMtRJ/C0RV9uGeumh2DEgfis4VPvW5TJzhLp2XEqR0IK2
ZapOUsr0cYKZfSUuzKodYwy0H/dl8d5iyCmEJRBgFVyLFga1RpVtuRMjKDeDQFbZSPvUTD3nQFM+
bwIoQmIgoEO1l5Lz5CvqM3vURB2Ddg8XcuE5Zv8QsGbVS9ZY72GODyqie7NIMwp9H8z5n/Rg6i43
pUM4PqKeWmSJGFBobpOHVsRvEZmNldE3StOPYpGc0XyPfEswQ0p955nXjPYYiggdnHot+0EWvY9G
AyvdT5AdT1C5hcBldBSCe6Vr9WPYUKoiFW/0OJurtupsl7yxZZVd2RtG7n2kR6qKp2X/b0sLYkeM
3ienFS7VeIbFJn/GwI/GKZc/YkdHkAlGOdwL8AJWfkg2d5i1Em7Ye/C3t/jsjY8JzRN0phpIaSNb
mPu72+AjfQeGcf0fieMA5f6bt2YD1arJXJJxDRGUyjQ5zr/YXLIqucfCcEf8shtMUfu3bk57qlrn
L7ydjb6334RmZNaLGaFs3FZcAsbB0Zht80LfhB0FVFzW84c9hZ1SxqpU1qcIbMQK1JpFMa35swGw
MRNBHQger4eMr5FDK3mSdlLoY1o0eznU4ixFAjZGu6UcgIxLiDUZqUO+a13QM0jI2sRCpN7/fXbr
Mk13oP7z3zAcAV+5v+J3wP4w1EwcKo0KMVGrsA3TaehaVPxc/uHVcjcI4N4QkkKkdy5jJPGojlym
i6jsfM1+4n1OeWy0t6Le9E4gm3SZWZHS88mYHXivNjXmkBVc95GU6oOA0BGZPUJJ1/oLqkAZEHFw
iZYut8KS/+YR1ydDwV0MBlLICh9gpuuJ2+sb/EbGoqeQGuA3gfG2sbHJh++tq4Z6n6aqi/XhgVYr
SDW9jePUyuX84Q822kwxx8JmovLbV6cBvFPkhC94hYcvNDL/2w2ZcTE8urLdTW85uC28ci5G3hlr
/H9WsqXJzVc9vQdl1LR62V0fQR5tX1tVCxAfCYsmigbRp+vvUjnc8Vt+oDoZN1NRM/GSEABNxGi7
XuNBZ592ztd5qqON9y8xj6ZP2GiAPNKBtEYXvqQdLxuqL4yA3C0h1U1TSCTiM+CtkvFH51Sykr4q
y0i8tvrxdj14WdpXAXC5zJPFhG8Siyh3WN790Zi3Sit+nrTRTYYFvasE/t6AZ57J5DRq7WK2iwCz
XyNqxLXlIWDMEHVoKlNIbhF5xRkAgcMtplhDK+2iQSOAJpfJnVdku2i2xOs78itXSrrPlQTOMywZ
TkP0U+lYvELC0KnQpvHeFGWjIZEIBMiM18iwCHlCtsmAHcUm0PUorTzIGvUnkt+OmaVZFw6A/j5K
vDxDiwGUFSfsag4Uew3dRxJTRXStOB6Z4UTxdbFwdtxvwVxyZk3Vb+TIBbgKoEaL08kUuIH1Vzzt
d2Qi8POLhNRantltgCJB5lsOyfQTU1DJTNWR0EgMikcmigcCwSXfLQ/Q0hxDWgw0YNoZ70Sxmdc7
o6aDuIS5oAwpV3U4VuPl/GyMqa8PbbMb+nTEsGg/758S9xMZRs3LOnUPae9wh4f/yLgn9dGNHNmv
4gYiQDtA0JKFAy3hPzg/JECXCWTBFBroN1my2FKMmzdcT/BGHBOkpUNGgSrmfyw/d01WruPZorIX
7/pOjWCMKgS7qn9c38lSAp+e3GM9eNrzw36fYwdCnN07ly9F2ykINW8+dbX0PPheykBH/Vu7Y3lR
4FBeZaXigJ9Fo2/d6hzmMjolui0a3RTB40mkYvc01IMJMiQSv/Hb9TMk/fU3rNL/qZjL3xp2+Qtl
Zj8PJhsa+7oXUaMiTMnv6UivZ+8/3/uzw5ceUSoTaMyJo7DytyMbinlLN819aEU6IgOWccORflsl
srfvF5Y74fuYG4cnr19hwX7+jWHa5sAg2eNsM1BLBIVT8QpRBexpQP/1uX9eAakgygVVHgyOV3Q1
BqBH6yVfkNDhZKTVgZGKzSdqldY0LqDmAF5dop+4194QSRXgL1IpzivHVekosqh3s3SgttCFoCaZ
DmqvESJRLYGwvIThh/TnBlGknoqt0WXVhh5f8uR7XCbm2q8N5FPwmuWTExa+9qpUxsxdd+h78LqS
XO6YWiQ+uOTGKcX9Q8AjHgBoiR5OuFiPwoJDiKIiBlLLuWN4OVylhfYc3X6HbE1lsGkKxqZMdOmc
BWxOsgW+psbcMyDEQ4ZHHROQVqLP3p0mNm+MWtTqRN7/1UA2Yw6nPhSZZ/6jCGohOuffFefE9hRr
MJUCarL4eY/RFDpyh5pCT5Uea0mWU5xZwLezi8jrLRd+YuLIrN2DJImCHQGcWN6H7YK3hEw96S/P
TeSlzLIaVb4sqfMgyjzjiNcH/EIfALvYoSlM18THvld7mxRDFXQRXZ8Nyde8diyqo4JdZjFPKGHW
yHlJHv3lfWJutu4f26/d4em6rzNglbDgm789dWpQS8do1H3cuxHL2bFiborvTRs864usoXghhuvg
b/kxX2Sazq41TWwkHIQHTDZVIWCWsyggpNR3Q/+IZFV+pxdm2z9X11FhFSUkc7XkSo3ajawouTk8
I2sb27ZhhtBc6DFSM/4QwbUTFXDm6ryjaICIbat/zwVSxtXwF8FqPwLH2yKXwxFTCHN5avblass6
+jsZ5RHft23BLSY39C8zfibTSYJeLo+40fPL7t3BW94mGrht0rR6wClv604hsODLE6LC/wIHCZkl
r8xTPztdJ679nfgx+YV+E96CGAjd0WVTqXyy7tCFiT6hF02YQiu20X++8NVz2JBCcYJZIapoPID0
iMY5qMvqrU4IRmwQLoBx2S1VleZBHP9tY/AmaYAxdr8TltHampTFF8CB25YBZICxXU+Xrguyfw9K
sviDBB/0MrLCt1V+oDFtKuE2AIoRK3A5Md7WjRP/JYf29+tvoB2mcEgceviBTCPT/v4m2rfTLcQ3
e8W/EDzksAYcEKbgSUOa7CjhP180kNqtctG7C/1iACFw5N3HNJiOZHxWInmKYRSCLxP0LKmXCT6d
n4SBltZdnmCV3siwTlW5M01dq9r2GlvFlpvQ7AQbra+BJ/2uv2XPb0tUcVTJE3EYKdmlPlxJlhYW
xDmDMAoT79u95G5P9f5ou3raIfh0LaLdv4pGMX/IpZWRdct0s5dJuhZBADTBXd0icxKw0qJG+/pV
Mft7OYibwwYVbtxxZ8DWqSLuVT+UbiS8TZ2I7Qf/Y1fqHqn8qKrVixRFC8bvhlhNvKH8v0WLlqCf
+jUoxY4cCMzBDRFuI6rm0ejZTf0g+5R7Yznr7/2j8BNC834ONwBU+I5cO4tr2uMIE8mFscXYe+dP
qSiGo6F3Q96w4OtHVoEflKmeZ0f3j73aLTA0PEJugXuQgU1L0joqj/bXoBTIxv8aN9T9+xSrNfgK
fEZqqfy1Z5c85LXjRvCtFTgUrdesLxSvuPH+5KshN/kU42WvPezsHaf9jVvKtj6lUFJNLnCYhYLG
GJnPudq7bySBEeACTK/urhqoTfAgSaB5dqQet+jryPjEclk29prh7BoTKCR5vOmeWjA+ehi95/nT
otkw6bWAsmZbszMz8eXdsMBNfa0jXbhzK8HNgyNn2CIZrXXIfumMLawZi5arog5NruAvyGfjXrEy
q9v+qh318oPi/00d8tIgMtDftB07RslaH1OCAEWcRm4O4LLy6sAAfzkZh8jWZd+sS8dh3tiukfgT
+6WulB/OUpMDyTuAil1jpehzIPLERoj3M/LeJYlXngs7o2CzxPeyokJR+1N0Ux6peumIZbAdJkV/
/KwCKZcYd9zae8zCC1zPN3n+4QaaEg5uYQxmKOm/M8RBKqjIJ6UJJ0cF8ECCyVxz3tLQtTEj7wxa
q089MABNUaOYt2vBA3OgOXFTbGHLbgw18AGuQGuWbW7wrZcHFu5UD2wcKxAwyN/V4tdfa/k1oX7l
GzV76igNCF7UXzHdhVlralFw8NZVsGWYWqBIfAQAmn/97g5himh03CHiwjw8lR2UJkaPn5IzKmjd
SR6OFofTSNQX7yEoM+nohk1cDsOeKIMAw+3pIfDLCtkCPuu0XkV+qyhP47rh6gxtyTYOFI+RuNTv
P0u9CVmAEau8biccrnQkzd+i2Io4Pdzp9NHaFX/E954V6e/uQfFkbDH70UNgvz+A1IR7TG7Dx+9n
8wbb+7/kFztb74FxeFoqH3iXVEgX9O2+cBUsDZG+GXpRRT1LvqZ1ae8OeJC8W16Egvu1Jltipmvo
C5u2jJvgH57t4tYnB98SrYrBLlR0T3YtitrmIWhrMgV6WaeWAAlDzy5VB2zmC63uZ4ct1EpNJE8f
j39E8qNdMnIA4pSIGQ/58T8t1MVfFX3hQj48U5GZ9pYUjigHo7TTXl+9GcsXE7WLW2c/7HuJzONu
FywF8tAWGS3d7U1Mmth7YfAEmveR3PwAzXt41jr7EdOXmAvFyEQJG+jPVwUc9cvVCcyeUBgxchxV
QeqianbE1m+nn9fJPVYhbWQMhEBJWLnwvdUnIEKZh6mmTSUCgKUH3DarPx7lOlCxRqeHPF+1S9rk
d+61qaoHmBSFMnWUBrcTZAHx4hD1ZMCnYl7gcBZt4twG3VVsU3j5AA4Xsn85H4E1AG8AE1HESJXQ
oOqxulNrsE0d/jBRtZb2Z7CXnEcT6GFAlKIbeOOP7RHZhKLvGJiWdLHmg9A8gJER7/hPGG7EiWhu
FfnD6Mwz5EF3KJwDl1BpMy/AQpgUtMlN5b/DcTa7YDWc0bykhOE5vJdmzfvB2P4G9vZQhF8jdzkt
yukOr9lkkXqeeKRHhfEy7ub9fqFo8ZFjdtuVwKECUlpOYUA5SxLNYYxvH7GBCnX9iXUbTolrbghr
BIx2v4EH+D09UP9Z3NvWwojRlCSXUWHz2IZVcsC8IP14a4Q1eSQv4rm7gqILZYufQdUE3b57lG8K
w4GwXYSHQ0KZB8rF5YIB0Bdftj1lgDDcIa7hlLb5QraiXQqU9aN5ufcIValZL8s2NQ79zQjD6vDA
kD9Ya5qa4/AQH6udWddjqbkiIEj7f/RVNT3qi5Y2DQq65Y4eMaN7Q3jCmZozeD3HTgu85IJr86lz
HdmE4oNdf5WjRe6G7ieAu3aMVPYRuDa89gKDHoF4EkZAr2Cdp1DJ+vZ0GdTLe3GbCr6TK47LMUIe
mFfBkFuS93ykmpfTGHOSNJ9CcPRQSJkvGFnGR4PmirOjSs8+PUzgy6mC87ENJ4ENjd3eLYb1MuF+
LUKxwd3NxvKJ2WKNvjtE0lvfWZLOPIp/j0j8rpn2+tFgR1mygS6NE+YSJsBmkSodv3bCuY4inkXP
zSCzn1duSCuiTAOwR2dtvDNuhIX996PVamSAA3j9nYN6DYZOzAq+fCSeeHABCIwcpGeEyZqinLtc
5Xdtl+HTCIHlNn9EqFT0mzkXycwpj7GW/4wkUGND7ish15mOS8ji1I6fFk3jF6iOfWckembG85WW
ii+O7mfUAkiCAfobmOJZVNlXsnV7wgXoc+k/s7PFyQ2+/Q/79ZCJwCYkWv+T8JKeAaoJcuPjBlFc
nqcx24TJBcPg3EJQkBAqKwMKymudXbCR4U9VNE1PgTwPM0QtOWyS+txaZKRtNtng8sgx2nuDwJ08
1Q706f3NRRJaAn9yMmBoYp7qWDkL1l9QDEBOrdx4InIpZJ5DeB0DHBqFsFYHI/4e0ZGO1Kw5QfI+
YbfD7PBtdVTYj/uMYluLvPXGf/TrRgRvBvwjPtIdM6wjr+rNQKIDf1SWxlzrRA6IXJT8qYx/PlZ8
s9Ko+9dkAOfPWTt86ZuPlvJcLM5mJNsQDxneYlaW0TxPSHjSBElk+1mXdTiZP+lDRrZzwvX1QoEZ
OMTARL/pF5TW56fXQWux/d1xBODnFz4GfIbINsJwlmaumz+UlxxgOUPPchVL+b4RiG4zCKicHY7C
PwI4IuWmYUyHTjzj6yvDjH4kA6puREO+sXTyjvr0v2uG7F3QDABVxy+9PNDOmVM5AubgHTwSFsSn
/6q6091WPCMwrc74sUhjjVWj7R0vW1awIigPFJDZTZ42wiR4O4Q+b8wDQ54Rosl3nF8VMCOu/+wP
9iFDU2AMS6bNLdrkZEAFAjThOP9Mnv1nwwLHsMiMpohl3pVahsaYRkqoKv6mMItVctMVKEVbwZnr
UwuMXWOe6XwW4G2RbQM4yEC1hKHkp97wBJYRhp0BeT+r8ilouzqhXH3djjLhxyi+DSV/5DldHiAl
/NqooXD9KxH4wPLHObmxM9u65nzvfEuOJQ70uwhJ74NbmBQWiJ3R6+4zLFBkwyqtfHFXRt7oLSsC
LZAfuGQqWAmrAUBUnWAwNbZ+MsWYklxyvsP9H9d69WBl69IKPXUSkgFeUkt3VU3XRU9Wrp11nfwn
gpZ2++/JfbH0BB3Tt3Zzq2D8pCjhJS587sMBSv7ORHFg9sjq9yGMq8B1qwPHEv3qKkNCOixltn+h
5ORUroiUzUeAK/8mpWzrEijXyQnFykF68GaAfoOwQrRjZ6A49FtWgX3i7nDLv8RQslHc9pU7QEcq
3nQL4nqNuFWLjtwmzeWmEJItPtxmM0bkl7AaXpiW2NMuSWecI9m+ZgWibf5lpS/pbQDTH75qK8fo
nmYIL/njTzTzHemEF1GryQKjCftQznLx1CCgrMwY1uIlYnK5Pnl8XSzfd5HnrLOapO+E4yv9ApqP
MaAcYBrmfjU3LtPfdjtArDkZm68dAPsd+qVo26v886O3yje7g3C12Nx6C95HTTqSuI8R8i6MaGvr
UzNbMmmaaQezphfGdwF3658tb//58GXPskMFB4N7sZGKvdqCDBE6kQTrSqWyYN+nJHVGX4zWyYXQ
2kdWoAStz1v9tZAlbcQjrFqCSgxXDjcJ448SO1EqbXSDNwvNkXqxaj2wFBwOPy9QHuEZl9LgeB1j
BCTCYgGYevFkRtWRjtBD9IcR9Fa3w5ZeCRfqJp7e9iM0xrGZ5tQtl8zElY67VsRmiZ0evAIGkToF
3V1gPICIXXTeyQvB+Xxpb3qxWBOCa2LfLf6uL/SiZyF6x6NjouiRmhyvc/bpparM1EndqtYtKHob
ZX8J53Z9OI/JEM/19BQCG0a+EpN/zkVtk81h/OLs/V68IoaZ7K6sCy8myknLAQUWvs87xCo2qO5B
jdmAF4dok541BO1pSvYEWNugZ9Ns9My8IEWM/eId9MJl9cecQC9bc2b1+W5OSN1o5DDo6K6/AIf4
B5lSzICSlliZfOQSakFvXRA907QOf1sUIXaStcvypKSSQW1ONbmrI6Cm2F7X9n8c5ZPBinEMZDN4
BklVHeyOogpTmG+c+58osXejo/oxKUBirS4mU9HZYvxlP1GT1YJJQulgJtPxcLYsdhOaR5H8oepU
1oO0vAjJqzlub0ZqDGaWJxvN39kzVoExtU6EpRquJzYbBN1oUiPZ66oQzU/dSC2O/UE8QFZhCzjV
FUSCnZ0SFvJ/+nIgXciXxywH+RhkXoKzMwaYplRnZ6o/O4nNpxnPJwQOOjDXzyUdmdmhPGlQTEWa
KlzKxPgHTl7kM4pom24WeUiECpAN+UQAqnitxMWutIZ5fEVaeEneOE7VqL0P1q5YgWQeiT/F4B6N
s3vTlpkFp6vwySIoIshFS9MD1kIQFjKg+9xqpmynl83c1axeEI0aEQsGZAgKiXsv+et/nTy0qOE/
oAXu9nnjwbp/02uL7nFw+ivwbkRfpvL7T5vYzoTrrKU5qOQmomAg5stxn25sz0jQxUP5SIDUSaNp
Dsl1BNH8p/gSKg8P9+Zhm2N6Xal3PWLf9pMpTeY4alZnUQdvHnlwEflPlpRAw52fHNewnNMwSsY7
afZ0c0G5zUun430zqemuDTwbubWLGf9aFon0rXYwbKbXg456xcPoivhgEdYwa7IHDJJk/SA3EOxH
awcnrTTdT7xVhtMurCtgQLr0safQ8sxXJY8hl45ldrOmBuAQLvNDu/c3VXB6mwwyWtcmwFx8rkB9
zCUEt8pylNFAONj4jCVosgA7baAOrln8bbDz/91ma1fN1aGu60IJgunTjQWbnRKYy0iCISK69sIh
OhukdeCGqG5zgS1CTmr5wGQWvvgt1PBJlmdHY6tY9xGa8gL2Vmmi5J6iQGV0NvNxUqPgE169wFBZ
17aG6DsMBN//6sztmxxHTblG09O0J8Oy3Pz2Wvd0RQxYnJ6ubfb798u8StRnSuC3satpA8HSpBvW
PLmz7ccx8X9bd2SlHfy5cYis1gdr4ngPcxWZh/W0mSHp6PQ/fMnhuXzLcubMb2/f5Qh7YLxTWFa8
qwNrVbLlSxdxcVri6YCqCyktpzOCjwq1mfkixM9CtU5ScV7akD4eLdgCMPt7gQnU9ZAcnV0USTh6
mcO7OOzEv+h3vQhW2Dj9CjjEop0fcBsWj3SxQN/myrzuMp8oxJEK13NH4d67l4ibqMI+Q8gL58qL
p4a3HVWIST9jKZMWjt1szalwJWtu7BuqTHPCQSVC6iXXN0k5QxSdUxxjUNVa10yCnmfGHy70rRal
mcp5+YfhXRB1SShZAOcoAvBB4m+iXwPW9sH++/5xL144tTKk1g6YNhq1Ehp3X/00F50aWzGOFm6J
cytSHlrqPDWMRJ/HWIeDjB/vneQPBuBiPFOHoRv8xO3BDo3OSZcyjx+DuPa7DqONfDCB8ZE2lvtx
TKqwRS5FFC2VGGQmoJ2qJSQGA3CeceEkIlyD9s8dfG2VmnlBj+m1Nt280PwUu5SHVX9nUkY6npUF
7TqWYHiaCjFF9ROqfXh9R6YfZDyJGW0FsRNxMY/lGwiDeDlsc9r6fjrKHAjXcmNZt4iI72MTRdz3
42dH0rrFlstivBgWfeoqU9Fwz7bxWma39u95Tp7XGiET/cqS9KZrhoUVR2hi7TgcayyVcbljRPGP
U2zNX/GNab4U3aI7NMNavAQ5dMvrkFT1Cw/x/0lYzSKDCrTSgZJp0MLRNI139sLCH8wL0CyykYKa
c47fQhfWD64zssmTmmUwZ7mM5j9pStPikcLipo9E7dtjlXHyStYiWI3XIxFO2jcxeKYPsKOIsQhJ
2dsnWe7NM0CmB5qqFkx2HulWe8mfiTacifZbfL6oCzRLl8mZbD6MyGPqu61yI8cHNzogU2N2qnRV
0N0ABCQhPbBFYjwXeKsn1/RCUfIFe1QGYxTg9CCAThVOhu8SHq4edL7p2xRCcRh7Hn24r8DOKXBF
FBkwGqWUJRv5ZIJVlCMWAwY+X+dv56NXORWjDkERG2kbpKGwFbKxLrxBatIO7NDCV2MbtvlRGbDS
YHawnXInUWHDnHXPRihxOKLeJUaPmM+L2jfiu6S+O72VnadO8IgJdxrjpqjKpYDxcVxai40Rk/qY
BuffvqGQG8mcLXLJkn4YuNO7RD3wmTczHQhHSq2OtBfcdBhE3GTgy0pMmPCWEderCGzWo74PoHBW
GBTB/To95Mc+jenOOihtGaNFgUm/JdbPa2xwlSnyoGTwYPL/1P3kRa3k8Dt4xozTMJgr2deKpiJp
rrQN5IUyWoBfc1shoAc41Clfhj56UvVjuoI4InSJ6K42amivDy7ni7YSABLgMN2QKoYsZFH0OjEW
Lz7yOpzFK2atpjXmmgk1F+IiHhz9ZoDtmFkyNtV8vKdBJnU+aKRd7a2u189HQk3K9+mrYjN+ktuw
aRiz+a5OSaCZfPv803SaaTaAiJIwYiEV7IUu4S+H4vtIYEyP6y3LW4LDabfA/sQv0+OEZIZARyJ/
/4IDXR+RY5EJJYI2XCtu1UdKQOGZeytvT++J7Ook82QcDDcs85XZqkvpmXQbPoDkv8RfGJGdMmkH
rT+IK/agKu83zddyjW+fcsJ8rPgptgyZWjOi6aJcITae+H5yNxllaXXUte7LOYu1hJ44m5KDLgPl
Zo1DlfnhtKGvJqD+Thi4w/AsSwuCvaSrK7xkz2X+5fkZT9CVWfUskPHOlJ7fFqepYiGrFU/i3OUV
vXyd+mYOTAnEXywiY7eFEgL/cX5wqcdIJD24gjGHTSPxxqXMr7dxB5PCPIsuWDLYyEXlcZR2kEUI
hCGqTYz+ps+avFPeaiE2ajF7gRlIZOu4kP4Ykhs+VMj7YRy/vWC/k1jB3fgqCxO2DKVRhInRQsgV
5/vqx6rG2EA6pHb/aUN3fUGJQ9z2VvQVPDpX3ipn4hF8SqwwNhe72MQ7xSi97paHyG+u8ZjofbMO
R5eFbCF20v4vAIQKglZ5hahXnbNCHsDLn2EZCdhUJdgwOnlNhs+2l0nrAhUtVD8zReBe+DZBSswB
0B/bkWt8jpvR4f5kIdMvVuhyY3JfutCod2JV8kPx9QSGV5zvlanJaM3O5ORg96nZZiq2hPjUt7SU
J3SDjLNieIjivYO6rG9b/7xdn2Ajze3DwuG1pcrhlyDICwo2CNVAeYQtKXssS3PmaUdL7T5XOd82
8S9pnWEhNNzfkCx4/k6vIJBzY/W4QHuko0bMIANuN9SGI9uiBi4+WAR7kjZs8B0JC7BzY0MfmPlp
qH7J/tzTRKMKcJrA1dWztf2t2X0VfJYzY8nAsKzKYriaK7L0Og4SYUEINlheFkbetFHALvHBr6gO
KVQ0djTIbCQQqJ62EESYngVaSi6d32p1aKGt961DVaziQuvutAW5RJLSEXXj9MlODvbiYjOLd3Nc
Bjy8eqVV0DCaRij/gSPhX0AUmUZdYUh9RzPSicqKWyfhhwwaAEBs0HL2CIF3E4IhKeaC7GIcCylN
MPhKryzCcFvi/6ilyQ28a62IHDFz4Mp0/lqSFI15ut3l17vV67qmT6SN4/+52woD07WQ9QXC9q+G
N0uxZmJzReHm4B5n7UFGVfX5mzW/Lz/pl80pATEZbGcTKy77do23KnTkrZ0NyrFxw2cD31TTJ+Ri
TDdaZzti/K7JpXF5+750AKv1VU0cQudZKd2G8joKRLlj5S/QrWnCPPtsh+FLi3dDX6TBIycay1Pn
/PP3ZVxhsydKbWAwEORAwFJECLgaTTMdQ0cxOV37jlwXHEJHxCOYA+c3iUdVAmuNxeX095CIS5GB
RMY5S4yRlOZWnbN8AyZhLQPGLji6GVFkaNK3LgeceEMLvAVRELqXk5HqYWnqp7wXj3LkbgoTCIy7
D50RxnXAXgacVFrD4WBZcrXaQJkY3cgmiTVchda/fNkUgbzfGrLh6ptaaSO7kOXXeJdPrPyfrklS
9APvVhkqniQ0J9taJ4E963x48fKWgqnI5vrDDbajx4UdPcfMf4sxW2fvCec5VgRE0y4n39WyX4sC
bAM7gq9p1jy2y1Oc2aBnA2enS1bU+Cjsyuzb790yHyqF3tOfkW3gWhnaDppaXkiE2/I6vEkkfqRK
LnruWtL4yGqrh2MxNSZOg9N0rLFFEVCKOGHyruOu05fY1wx+jrCzFRhQr1b5hV5SPipK85It1E31
4CY89+eN4CMzeANHU5NIURk/UT8qaJfU/s+t74oIDPN80XTdNspZKHJmEI7g7HeQnSgxGhLRwNEZ
H57GR5NxVLBU2C8M5d5ZNEsJsjywxj042rgazM2cNeI4piXYK20TsnLaT3fVrB2LISnhUHKrPoYM
yZRJilFmVNSzPNjnEElXu82uj+FfKndqnPudW46a8lh8XQWCnHTiDDCkCxuRFVYn0bGAYK1FkIum
5wCMCKZCY1Q1UHZKZxjRS+MLaZK83pWfTL2gmjKKvsM5RqHLxhFXEBO6RBF+gdEeWGtdURKZW8dz
BErDQnHAgCGaOu0lk8lvGcJUKGiY20+sjRkySjebu6EgTnaadpu8cbJsVecDGnvtkYWZmcuSOD3t
s6h4bNSA/mQgZTYo7v/CRGcSVMFbGN3m+DqKB+GAcUTDQDG6Y+LrXJPhiFr5xzQltgSamYlYXG2g
GxvvtustRmaPJz96VyBIE3F2EfMS3g2o4APGq+h1w/KaXxv1gdbf5BM1FzmZB9ZOLnY7Q54dSpr6
TU34PFe0VmCPJNEJJ00TZs1XPqCPGO7fMpllmXB5ikQZgMYZWNfYCLHqETKof3+MLAE9VeVuhFOr
axELwgoMX17q1UKYJkFp52ZLKwGlE1iy3eZFh661BG97eED/rBUMr8kt2YfrKFd2oQwFi0CHGLjj
7fcpUZwJMo/IaP/uwKecEjhFcsHJZxJU8FI6alVWWJjyzCGN9s5EvAqgrzRi4W5gel8zoU8IvdCl
FE6gO+OsE7f4cWUSrF7QxDlNW1+7diU/t4IAGkNc+Ilg7Xbho4cvfMSHDZuC8vnP91w+K4IOD216
SeCfNcZyRUnlWp8YZdiqgfLXXZlnc/S7c41zBwd0ehnci5EmL/KeEZDpAoGAEJSfAF3p3fhLWvex
vUiZ07iGyQ+q9DClnodcmxs3UN0fD3wDz9esULRyZSKoXTkt2m8HTFlsyqmT1eJXHlwQjaO19PlH
ZtyYFe1wi3IcjI/g5BMLm0eUqEO3DFcppU3WOpGxq/kirtIqbCu0m36zDHBBLPwuQz/4CGFai4uq
1cGnSJtcnOvH8G44tSAPXSKYhBjnxv3YWoIZLjVPx2u2wsbBTr33x5vQ0cUlZEBZEs+aRXzk40Jc
jDuFgqhcHzsqLxusDu36XwfRJzAnjVVxx6uB8nLWhThMat6cyQwTmUdyQb48K1QL1Li85rtuY/yM
Sm17S5pmw/bdZvMr5P10aX4d3y1gMoRjAajRNmcntUY9ow/fc+dyvzXQzoZf4aga8jTSYTPNA5v1
2/CEH1+teXVasvm2yRPpEnlKPCldMcap5Mt3YVcwZuEqtt0mI5JkogeC6e5YScmOcVsm9z4ITAef
v88MvU1/g7rgiXdkQUGIEUp8NsNVH0Y2ksbCsC9rJ0H82m+CC+5Rf0vB8D/F9EAIeqs3a2gJsiBn
HTD/i41zTFWKNw3lObyH6u6WD+w+c/H0GZpQKd9TwKUyye226NVEYc4SG3eN9oG4Qbe1ypDJ7n5Q
mbL1NkJppulokOlt0Gxjcvuzb5rBdNG9Na1VAYYahFX0NL2Pj+UWGMPr6o59FxB9zrOgtphvgCqX
hNAC+u+cRocIXpPt5dl0dAR3fMc82gVQcA8t9AiKM1r7Ix9pD/2o57HwfWOdE8WQsLu8dbYzuTOh
s9tIXQBNf9qkkdpMzMVsel/Gcv7mzW6xFYUSsG/K1xwdk/D198p8MUHO221NIJJp2q+4buCdVEUm
H9P/MTXsin7SXfgrCFglEZJd30ZMtK53U28OPW19t2Kt4UAITZaejVkJvua73woZDueMA85EPR2d
NI+4Xb8uGhc3pUcKlxDiSPxIyzKsAzBZCb5e/sTa7Wza68227M/7+iXIfG4mH/OfaYnfIRv0zXgS
dsHn3cWCKyKkcXUqNsxnNRRBKr4iwLdSjF5zvVhVR6NX2KToWwjKyJJJX133ew+yXRxkeZhLjN34
X6ybzBDHjw0bAeDiH2ZnIfbo7Yp9jh79xHJ2/BorU+rmnadXtCECmoiShN0W3y3vrH6PwPzbBWdY
pFgMT3xZmZlmNVvhge1KS/Pu6hqF3UsUu/21Ok9vG/E0TK4ghis5AI8rsF+wH9GwLOjMaVfAm2j4
VrMilFth8+dEoTRURM2u+1GoGYaBHk/TJauePE4+ERLcS9HjA1HyIni2xxkWiDwMLUMIsACV+nYN
kLiIBjywRaB6p+ZTupCxOz1xW8ryibH+H27hwDz+u4xH6vGeRqIzYns9qzR00xOM891kUrZBcZop
349rGG45HnXMdG4QUqDnwfPbiwvun0KWyCB/zrHhMSoW9lUYbjYOFV2zH+MaURdu3qm3w9A/a1/R
FZdqLjNefdWhqc6a1/2lZ4BBsYHvnJ3fkmgenS+Cs0LRFsX7yg+HgHACMR0M9aEwgnJILqIkWtNi
EPXnM+MKYbEaOHxodUwrZVw+bLG2KWHafULAd790/1UzTkIhL4IqzdPCVxtaJxvn8rtbshuxTg1D
IDk0YPo+TGjqvMfxUBVHjn+PpWx9xhrKQxwtiZpcGVlmqAKC5M335BL+Bp5U/UUtJCWJM3RKUBe0
JA9nMRqT6xyllabvC73vfEQvR6JlznTw9G1SRf9v0dpL2aLNydVYnAInG+SIRk5bZZIMImNnLVmt
ENeFJ+rsEMvfoNAA5Y0/0tD3Lr8kXAP0GBY4H6m97i7Ir3b0b31fmYSRJAnj14svf3lHcqf9I/TK
cOGD7Q6s7N8QSmllmFO1tVV8N3cARUd+70s+mJ3tH5iZ0DQsfiepK83Uu0B9VZVXT7zCilTlL1di
3a63fFbHmKfhPrCBuH6lUZipNn9CfpBqZrfFSiZRXlpHZYunEl1TnQH1ZCUUN/BdeS/fQlV17Lug
0jBClZHvDkLOIC3QprxT8d2e/i8wVzW1YbHZ8B//+P0YYbasdFPhbwI8FK9WT+PI5IDI/C1+S2VE
04jaDJtK7zWVlTEu/bAK1Svc9fwB0lKdFzvoxhWULf3oNya9hCfObL94G9ZbzVSMAH24f7khDRJD
L3DQAZaIMktQLfF3DPjSAG79COwlelVlREChsyFlIH5H8C6VWlAJUh4begNUcRakAYX3xvMv13wa
5FNil1QuF67oHIUvYyIhPu2v8tAqUbYhWGJyGa+8r7zv7H2RV7fi6xr15zTxV26lGklZT4xLoQc3
dnfFayTVB/bft8Du9fGFif3F+NcidhInGR2ANAId6k5+7V0PgdKQrF1f0ALLB47vb8xMMSaV0ZDs
ZioUbzpSPY/53qtLWC136SNIijYrfFNis11ipTSbw1c4NhmzIaMuERPnS1Nu7F/Nv8MiPS+g+lGW
slnAnjos3lR8+SsJuPZka3/WPTkjYbfUOjxK3yULNrupqZJALWOrbR95ZodaYxRya/SH/ivXEId8
3RSN1C9i8NHMaqISLIWVNS1eXJ0Sf6nGcMw5zXwVXjfqlWBfr+J9FbVzMx9aLTaUn1aL/Wbhedmm
d7LUm2JUECCOQOgYROUKRCvSADjD+vCHBUcM4bSWMcWA9HmPx1b9dER2fpqwQwSY4E6K9b3OkVQu
G7Gdo4JLd0uYQOI3Fz8pxpbj+SE7XCEud6Tq3robM6ycH1rFS+1vf8La9UHsAeOVZqO6c8QCxX9S
62SQKOKeG/WHt+BOAgc5PBCeffZVHsCVz+HooabYPRxFRT4juUR4OBvoTRjFs4Za1hd1vB0uSS2i
nBKRhf/P6yo9isdav/CP4oonWeCh7vIpMq1+Hb3KDr3ReilVhevQo+i75XFRbQiy+3E0ZShZufey
lXaM3+jaHijIorbxRSDt1cm5OtHk/BLkoW/V7zGQbguK8NcvyDSzHviv/PD8qHmCIdV+NMlBlGc3
7dyXyqYCHQt8/3J/Fm1+fI42eOugbJ0Z6zli6/F4+JPrL84IY/fRbRpK9iJqxIgpG0aJhjkndbHh
BzeD8HsLcP+GPkfZZ7K+o35D0M7Cy0ghcG0OFeprVTstLTz/XetQTgmppPqOBa/eOEE6BR7/7Hmz
F1B3W77+Ij4X+vPbWHCeub+ron1Dv/ZojvFGOm6BWRwGNeAIHDzSN9Uvle+kVxTfFJ2Y6bp1VfU+
YlF1bj3zPTKNEFydPrHHpWEeGSy0ZLTBrC5mGEMRfRDVNqN/DHYFL5DckLmx9JZmlzNLQUql0/sT
hBiPX9N3moBd5xINM0C0d5U/6Ek9hyRprMdSKx22Lwm9aEo8lf5Qbi/Ul1yUc94LxJes/4UE17K/
5wSz0+DI6SHj4T8dbzN+LrkjsCVR25Pe4uh3kVJWyrhhLgJdp4ljRX0IfT2hsiknh77YdPKWCK8a
+SCkW696zqs/ig9xDK+Ney+3J/4/qSmzuH4FdIcF9QD94W2avcLypMYJyzF8iwGaFs7C1SyjFpsu
AFTlj/o6YurgP4Y37uDpLC7V7QsBEwECddhe8j8kLNAKbS5dE94hzqjSmGjGt2zkfYPxzqvTuo6X
kPapryxF1LCD6G6GYAek+/6K/k7s7FE1A9J8YsgS4VBmn7GWdcp3QAyUJxNgw2eBBG7lVClf7WBW
uW+UAZZLUsz4ME9WvgS8vak1ihzEd6rfq7txQrYS5PeJyxE8kMFD5RKMdJEXnslpT8xgLw8gUnp/
KMVtJGbTASAX0wjd5THgrk6xvMooGtZE2EQ/XZeskWhXoFlPiaePykXeDfzMJ1rJe9IMv/LrN4or
8Aq/DOBMTgjEJdfWuKJEzk/rA1pqJm0sFM9XRCdIsGRBGTAds2Dj5Z+wWvrcjIbor3vVn5p+Emuk
YFfR7+eF886wUKNLOlXmpptdrIFLW8jybkSu57GU/qMbWsA/OkXGmOKr7SoIIdSZa7nJW/RicICN
4YBa3dQOTZDZbcXl7IZqmDzXI8R4aYcc9lChGvq7MyeYscd9T4e271sqF6ejAhqZ3wcS3Q4tylNn
UaT+69VMa0csnVqsYqo1veYWdE2bgyV11cX1Ss0IwyatpNqdpIw0i9SlGNwghQ2u+I7jcNeRXmPD
sOI53s04tNn5iydeVVxpSKYJSr0UioLNepwNNAy/T0HEfyL2L/erq/OlxK7gr/NtAa7CXIshOCHi
L5KUsfEyn91OCas1FsXiLyX6ZnmaWLJ7w9ur8DxUCq7kk+c/1ptYJgc15zT+24Q/ne9gjcjYJ62+
vtaFCUJL1oWQRyr/gJLk/6Hx5jI6eGU1j7NtUCDKGZzQTPmDEKqYRrS9UXZjQ7+BAqnfw/ToIcEw
mlYriu7/+nFY8pbAkgku+sTo+pqLDaX2NB1+NtJgDtBmEp6VQkJU5ipWo15bdoE0qOPp6pbK0LYb
pocIMLwS01ZjtFRq+BoUcQW/SMMwXArmXp02b4qKeZzHMGUdA6vLe4FzXTjAQmTTFrvkD6ZUlSS2
lc5QvqlMZ06PvncYTyY5kBVIT10XJX0X4RXSUFF85fOK77brEJMK4PhlQze3YdshhtCdvxtAlfG8
YW7qWHItQXTqtHnbdmDQAUI4j7JLMIL0yzO9S6JDJX8IJcpp2SVEYgCPWcGWGfLeqE8wXhVWjOzs
1Yn+fNGOv+konGcv4XSPO66WaNf8Q21Echyw7yOPSjI7KpyEA3FX5V4VH6owIXliJDfKx0hD1DAB
Pg1dBCamvFUjXHUBYAUEqvfEIIckI48t+F5SHrA+9f7RWQnrO1WPSWPN9UcSvK36BBnxi39B2Ns2
XTt04oR+INC5uN2J+07oRpGwJ8HrcnUuGuYfBPtic52X1lS08DJUg+T2NGXHDZfcq5rm4RVWNP1E
YutzqhlFrP0b/aXtbiQINV6Pnxi3WdKdnAlyHpVsm7dMjmKKAjV1OpWSgeXis3F1dqnFi5H9foLc
vq+I42X2IfVIVvAjHTAkU5ai9iCWkCTvCrDni23vS6h0q+K4bHHr1MdB47CTUNTHNXjvzFaK8rCa
k6iZMho4Ofs2KeIL3G03pKejuw4tax3PLHTI5AzUSGEblBCG4ORO1cGnNcmloRraF6u0nC4RSdkW
MKDHATVEX8jl8ddToioKj9/rJo+tSZSuavjxiAEQbj7XaouuDUeBhmY1y+CQ4NOyA0cBOFgFS+ot
nAPG/2/0M8apID3nFdhYNU42iHvtDkqt7IeRzbcp/mxaWkULzVolaqL9xF+xDEt/18I598I+rtLZ
u+Uyp8aG5GLYBSouOy6FSuv8ykZ1hpRhB+g4+EtonP0u8EOSH6RozJg7VyYQ9fnygBiB3WdPkLRz
r8Lc350iKq7NY41ho4ROfPjuzQaOIXvujQjrMZthNL2YWqPcqOGaB2i6kp7Q17n7HyYfZZbtwopd
X1/RfIkexCqS1b24jfzyIOZtkloky/oeEOFFplZEwLojiwfzOV5Oaxr/Tlp2QVS4lSADPxR8QHad
cCRICreOc33lVfAHVvYQfuSaxtxYQFdfyJwIeWyu21lTg3WU605q49yyUK5kc2zKwSlCsZsTpz3l
ytntpOLl1jB5uq69TNw0H/ZT89ehBrW0qJD1WZqcxMIlcf6yaAVMhCfbLz2DbJyFVlx/aUFikYOd
B58W5A7+EUz/K+zXoJ9QMHpYY3JFsrfYB0JIC1SekA46HMLTW/aU111DWzB2SrfNGzNMi8Eh0mtF
JkM32U62CKkAoKrSChCWGV12D+4SxrOP+aevsOCO1JwlpbnFvJXVz6k972WLdTkcNWMPlxUb5Ez3
vo4l2fE7LOMtVupErl29yEIeGxqyBnsGSj6DCmaEDLOTN3jLIbQnFKEpSXvygpmXzBO25Ao519RE
KEjzFNn+NuiaVvyFuhwro2nImcco1CteNV3ybV2H9Uu9iYGGnhWWI7Ntnb7RsMldJrth16lUeYa4
g7H+T4PncOdsQoDr+DJR3vc01/ESBQaElrEVAIwCqx5vkjXf/2Jn9Zx+JfC+wcu3GbV/sSvW2KMV
jDsc1K46xSczBl05hA9V33KpT+RQ4KZdNpafZHgsY8XSVvhjpRY4nKmdJZ7Lj3mTXYEsiDj6pkZn
j0aEiRMZoBQwFyr4/XfDiVwH8siMgq3VNPuEVXNPctW4hK6dfCgNHVp/rinwredK4RAwUxNFys0r
uaB6CbbDmk+8WanCbT0+p/T9O/Y/zdeeUCHMfyfh9oMykOJpQSgUoNut0vEr9efSOBQNPrPwkOjy
dk857MiChpx1G6lys1M4dhYxgM1+TQIjAmxf3QSZtDHuoxHxijnS7CWcEc+CHZlkdTmAI9SorpE7
nekDnfEydwCcsxWjwNEY6J9bHFxIy6Gk9kfuo4XFr1ZSvYiywHU6c2p+G92uZ379wqv8Y1Dx5yHD
FU8yRut6R1lnnRqXPl1bkTZbxGXVnGM8m23BTb9bAwjrnBkxVDB/SeeCcXivhKIotiEU6a+tfhji
xRhDBkGUXYTli+McaLga5cXtEHUXQ+BqzhicxphUNRfunDXz+58MBI+/1wgBTQE4YZRIcqJhWWRK
oc6y1GYnsRG0aU5QkNvsrB1uYt3LEew5lirnDlqH2PwTReluPmeEVd6VpDluva/XNkl7oUmHckTi
+aBpZePcbhJC1lbkMx6TLMnUAKDXshthnfKs91WZll+jT2kAPUPz+De3Jg1pztnaEcI61EKcSHiN
rB9QcFRCV9ZN+zaUVX+Po9SX/Oma4bibsxsDuP/63dviu4spbbjHoN1gtkN9WaqNUruo8+AVbkdO
dA25QgkgiLOOQThUyhlWYXBBL0xQkZ/Wo0BPyrXs7vYawUOEglUTLHzo32gx/Mv1kmafTLFnSo5t
Ed9TyLi5Pfbgy6fAYAcGIFN4929h4oK010GU6tttdkE25AGqpn93i4m2K0sPDjVHSkTLRMg0Bdh0
tDFbPmHdYjOkNOqqSTKADD0EdbJdSJG2O4x5yWYeErOQXkU2uytjp1BtPR6QuWq+MJYNm6aXAMxd
R9iTDSpxkNrMS+zm5ZL5j6ktxPxa6EsIDveTKCaa1LYBkFrO+vNa/ZHPiMFibNUxSu4XF6x9dVlw
n530BCM636i5+i8LVSXnAtKaweJmQ9WqdAFBSTzhgnKK66md/cHdBunpuymOR8XO8FnztIS5oFHb
zZM4BBOggTKC63jjT1n9L4HAqTNsaiEVJgz1b3aVtn3044xeXBHG/mtsuCmeoATwh1L3zh/kUofj
LISeoHR72DSqt2YQkApW84+uIHcEtcNHf9AWUCRR+HhwE2bzDqBaNO5Zh+h67CfJtmjrMLm3FIgh
DZAAZK19NELXrvIkzwzIz6WznkE/d3DoYbZhi0f4mi4cnGyfIrpZ6XYMZcoO5qznZnnbbX7PTQKS
gIiMQF2k2FtlHRpV+DbYKbNK4Kl08359ETlWANAfSrHoosfYZk3e72wDVwcLIGNs93k+pLd9kMxb
hnftlko2E0bNOXpwVMdMOmyYqzZatu1MbIfDfAM4vneqqqeRC94yrBKF3jl3GANQTOHx1hhePd7A
+yMr7oYPDm5nn0L+J684aqUoaXNCxz7DYpgIKli/DU9czyaz3sQ5R3L7z0k58z5ioWDcqDdTuQV+
jXPAMvZKu0TMwaea4DYl7TJ+xLhHf6qsjPYZxNF7i6J8c0qYZOOxIMI8eUK11wOOTM7qRM1Diuk4
RYJdqODz3LrcJKi1IeLaYRePQy9Bn1YlVwWQ1wOpSxtZD7yRabxMwIvougGyaUc1urUVi9eZib4T
k1oMZXpkaL+BKOQEJ5CO+42KFIKnmsp4I8sAZ4Iim9G9Ck1lDz978lWnEhS9xe7et++CWML7ihow
VUlTsZSgUC82TfBbQTOnxVLL4iZ6cGAWgl6OjBK7R6jdb7NqSvKc8rQLmIbpPvB9BaBXOn42Y8up
SOkWe/+iF4Kgo8AwNsUvhzhXZc86oRXXxB9zj5O30JqJ9EQNWNaf+3g63pu60MgceLNZcMD8RbwA
/aHSHbipdJuYC7/uMhnzLR+/EvpDnwj+NYMYCWESB6t8TDFCwcdGu3hHwDO3eoN3b4D58RNgnqSS
5VLtSa/8CjSmKnqecsOZcou8k+XRSBzl5JnWLsujMlq6vu2dh3kY8IGeoCNak3z9mM/c4/Hz5HUF
z014OFhpUDKSlLkCaz7ns5B4oDxTkMtGMUVp/F60nROVh/SHiC66EWlJGL6/ThHcDKtl8iLVMmG+
llykDd7o3rWA54yaa7wumZcZ7OMQYJUlcuRfPU0M4tr6+YlxrmSiZ30QSTFencmFCsbx9wGzR5Dp
lH+UC1hvMIi0kesX3PVgP4VVeS8F3wIaJzNiaIEo6XvOnTCTj0mD/PZcH4e6JYBZVulyvhq1/9Gb
q6nq8ndvBH4NUhR/FDVowdazKvqpbKyIdFKheV+f1295q3Be4rskTNTs4prn89rjmfIvhQqp3VjJ
AdfOMV5Z+lk49Do1+c3QGtcW9XyXjv+4Ztz9H1fbuFo8tUjqHTggKwUJfRqZTXqeR4X2132G2BEN
TFtmLnFwTz5kPh4DpSZhAOQR58i0Gxr4SxT6ukC7aDVXVc/u2qPzA7riK/FvEpmqEFVMf95kAld3
W952JLl/WPjFhII4H+oBbliX5k1bvE84iNgiMbGskBMEy0Y6VLlL8U0zoh9YtQPbqEv5+ZRk/gMM
eBWEJN8QnJ+aWOIbS3/0qlYdh4GjoPS0kquAT5zfRHk/ItxuuytrjAsTpMUxIVWfa5abA8A9BJzT
VE/miJeybLSVq++ncheeVWvLVEkIj8dvH41yZhaqmfzKsDDgmZXTP4rIfpmUiiHRPxqaoPo9/oCU
Iv6bpLA1QQJSnhcXR7ih4qQrAMHgefSVNW7Vu0JbhodYy1sGEQfGdHwEA/e9uKiF9Y798wYP+0Gf
alyAVdWsKU8k4gGFh0fbFRMaqcO2DFIr5cosv0yGVgKJpIywnMN5J5I+K4oy0Azza9UOOcXA+Ls/
VFpmYLULNtBfMFjD4+FjnkOLZxgCphUICV07eMcNKQPLMKcbaQmnHgI7Y93v347zAk5XAc/rKhrh
Tua3cwL2cPaEhusqyhqsypqyPuBAN7WpWYClrP9QRVcoKD6CkqFde5pFFxKz83wMDRoW4F1BJR0p
7GhYwKIQ1Hh2oWAWFJ41OCn0yCX+aniHVA/MHbpsPknmNh6hSymyGaulqBrD7N0yh72MhAcKGbNN
dq5HEY6X7Evl7lrjJMm9Lj1iQUFto2tCLiKm4mHDQM5YLPUwOxrlLgwiJktMXR953ulhMfw4M4Ib
070vrTw7yVXyEpbKUxOTM9BbcbRRxTOhLbS/mqFaX8JnzI+osPJhuyO4++FJgZuci0Cqtrs9JtoE
O2s8OQr2FHr7LzAUc7gO2zv7BJ3C7oYm7jeZqC0lbVHjTa7wLAsoZlBoQQMcG7xeL5ZAEJvIUviC
jgah3yyamz0IMV1/+vq/bswwiffHQIJVxTzEDzWQD05JUNLD4/QpNONJNhs6D6ib4NHC0xRfNLmP
6r7fRG5Y+NOjIZye4tCzUZ9ZteyiPYFaY1y+SM19GqpHBAqnss8mkbOj5u60CkdYmvmhYVJc5F/C
wbDExM6DLT6t88+Z5yIze+fZkOgyhkEnc4nywXv9PDzYrrMbqunYIZbmw2dOJp+I7ykbitrbigTQ
rBzvpILV0Kkk+LZ5pNZj4TQ6hc6wdq2M5s4LnctVyuNa7SXp9/TK7yYzXaSNryC1Kcjm15uNx7Kv
G4o2f9Kqq0HPN+c6VN5y/VjzAEU2SHZMx4yj6NpcrxG4j+Xi3ZvO5IiPkzCbVPOjBTnMmSEPiuiZ
qptU8pwRDN9DbQr94+0RXgP8KmSY0l3r1l8iWq7jpvX6t33bbCKajNTB4ySYk0vmYzDvO3pis5Bl
OoJFLBxByh81EwM8GcM8vA5NhhQLjlkq1VtxzP1/FaORR1KNQv45rxEbM477k1564Zslfh6Gtk+G
SvOfyj9bgg3wY8tgLWFcKhskdsQlSkpYDBnIu6HnGrp41NLHgrwshIbAfi23Uv5u8xUNBI4AWuyD
e2J2OTo0v/tOxKrDb4Mc/SR6icl06do/h8aylSc6eMP41Ira2CMf65E86BG+2qGusFL9Z93mALZW
io6ai80pzw+v8WnBZF2o8V06+1isY2yAcLKh/d1elOaS6BfZA8Xk+Yar6XuukqtEGYPKG3Er54wZ
Pbxg+vnSmJ3JdQaF7bNSXYo+u05h6BX1jIaTVM3nqQwP7LQreHbHCpZBPR6i7qy0GMx/RVTQvzlr
e6+C+hFduJxMn0J2I4DC7b1Y9vqpbASmS24HU0+lN/XuWojYIvCTVjKdXrQ7k8zbN13EnM/UVjM0
f2Pk9hW4Gm9AMFOgzzKGto6pCI8ssD+IMF6Jukd0JlICz6w6LSG3tfGZXGD4AYCiXSX/p5X8+4K4
PxyUF72WUtdJ/LWHYR1tq1uW+6RUismIQ3MImSJUyIuUO/NYcM1woSalqzNik8cIi031CnUhcAvx
r1C3o3UzyqFnXjN2dQX0oDi0QAli2PDVtwSBVBjLfzQuRbwTQoWH/ZWCY7nXAvy/Z82taPGXgMu6
0svDa7iX9IvwjCqcTr25LgAj1Lb2Y/UazL2PUcat4/hnb1xlftdYSQ45s0fDzwUspOh50qcvTaWm
oVGDQwJLlJzpoRQZUFnUceAgMKGr0CQSiRoS2dXq65gEcqbnsZT+e2kqQGzT2QXIpGxUN35UYTCZ
Kp0NbYLeX11F8CIEZgjLeXSYtzf7zyfHJdgFn4eS3IQ5M2Y2s/phfKcYGD3olhwY5eMqGty4RB/Z
AebFz4wy9DzRYNhWjfaw8urZYgiMBcGG7ruFAKYL3dpbVK8u2x4RS/WpeC7kktfFleznUJ9qhdyP
j52pJColitjyquuWgJSo1bCsQt56behQ/kJlaZTnq+oLcOn5Dl8n/MvxW6vpnpGFcqMDzExdrm0G
JWQgZM4Bv1TUHwTqidwJPHsyTdVol+K9QaRwKBH1bnGpCg6JVewJhsGMG7MSow3Gn5vcwFQtx0lk
npf52GBmnMBiR5AYlrpeWPPdjm2njEx6DiqDRqsDV9NzB0HRWd6FZcQx2aaE7HULQjQTzinXBAf4
+bXmFB8BjPscH/MlyhwqvFf1PHn+r4Z/4C63EKeb2/jk0zF7EhmJ7qWdeg0ONIrZxbE2zquai+r6
ITygi2HahCdSm52UdqUgZNKTaHPbE73h6Ck4arJe/IRzVt+AXM2fgzXMGnHlOQPRFSUyK5yskz9d
DZfJQyewYi2ewsBnpJ+vdRvLn7QJtAYCSyF4SMQ41qrpUQXn9NIRRbPpr5oLReOjLmflmXQeeSr2
A8FHsn7GDSa2t6RH7Qo4FlRejLy8MeJt0GKVmS1AkTqgOtJ7iBDippsslX3CfAGrXwIhwSLStI6E
GCE2/foBXs5t6edhymuIYjqbyRqVjpx7osBk2pQDQO7vNyIYbI+cc8EXDy6YN/TIFcCdMQR3GFw+
OTTbgchuTSBDnVXdwOMU1u8QY416IG9DtUIvGkrQ2mogXX3ZwmQi6Zx9xO47grX3hHnNKUxR94ha
F/0IEmjSN/gWmUlnGL+/5/Fhgb4ASso7qiKkSFdt6bmGZHltorGIs9A1ZfTG8aPCULIo0GKVfEnE
9/iW2KmBNeJuZOIrlSFMyGoVDVZMMCNBSKFFE7PFRJAsmMqF7sDMhPMKaSprcNqkxIa2UeQPdNqV
+4r9hl40OHP6/mvWI/w6+DwsU+ioKqgmNEEMufiYan5huvY1c8ILXi3Q/0g3BUPE7Nq92cTzIesg
RpmpEr5L+agk43GjY2nN/ZdLfebX0suLu05ABgf0akJ/u6z40/zStfoJP1HLelBBE7U+LR2tgmd7
hkSVw9Y7pHJyouzZme1v/8AgmPYk/8oAoE/84Gn4e5B5OUiQ8uMlfhG5BuZliPHm75faTcqbZNu1
YaPZqoXJZ6NeTAdOnKJTmZuh5RAilJ/tAtJ3ddh+/Bc5SbZ83Jvpap0+Tr/JYUGIAxpAo44OcSRz
LboUN82QwMPRcPWrdui3Kf+vHy7E4rk4uxMcyEAuYpslk0koxL9U2csMvShYQdM/f05SVDR3dmL/
Ny5jknp5zDVB69iv3vn0V1wKiI6bkFFCyqW6DkxnxrqtD/psSkOchaflT1t3xKjcPQitJj1Pkk2Y
8/3rsokBzLVzX0heodRduyRo34rqFVyMErVqk9uJrGmOlRNT03B6XrAChvG1qivh0nbyUhAJyU3P
sm9BzVq+7Cl2whyCoOYnaO83AWNgnNRghSVVPh1mX8XdNrdYRqjq7NAkpl7Mmi3tKzI645GD0FdQ
h8CbOqra1YkOgYTO+aFh6N/zXcua3Ym/9+dQ4NnYkihcedlmtJvGm7EzsOw0+Ip6M5EgZvlimvCI
ER10evAyQ1u65vmm9laosDpU2EDGCkcHqMLrSsh9CGQkVgZRHn9gJYCPiNY9gcaR6rTU3Lvc7PWP
ssgqh8Zl7ggrabWKd7r/5RQt8+daAtXCcvRI9lHzWd3aaYa6O76k8WRGdtyEk5Ne7Mgolldkldf6
N3J7spIpWcilry9YMZonARgWZSVgeQAxZBOco9GmxbYFoP5A142UWqSkpm8KAGjKs3MOxVS5lcms
X60Ohbh/2kzeoMDJZeju5aThG91SD3GS3YAoscexlBlTTcXn8RX1uePz6PxnBphXEYc3ztv+4Ec0
Kuep5edFfvzm+qD6pfmHN+pft+P+LKULCGLG4w99FZfWIJNuvV/FI4maUrJWQsS9j7Iu9lEzsMds
k3slvmX2993NDGsN0z7GQAh0Gdro6aG4aWhZJZJK9+6uDLoZf4Kgoj6wdeGbwMlRYWObas7K/9Hm
zKBLwaxD9Uuifl5A6hnjEx9KhHRSEnQXBaT78aUVgpuh32B1u0GfMm6qyNSWHj7KZSivfBH9UpF7
5ergFvzDVYVpJ9gJxz9A3zA8NHuJhokO0alKVVOFtfVDabC18/frhEb6bOrJo8zfY1H0+dliCRqU
o9jg/MvEYcSXNqV5Q/eiHNEu9rnTTkQ3VyN+h2Qq2rNFGVpYRRFbnYOMxzGvIIuQy4RC97cErDoa
PCo9QYqLrY7v6wa/3szddBLZWfVl9Sn3sezRv0dL7KSbM/oAtJIiV5WfUwS2IEhy8kufIM0/0q0I
Q1ZR4kXANwmSD/v/y1UQ5KiQ/TmnaZwRD/NRhuH8fY+fGJSakR7DvqesvSWYOljacYWACWiU344x
HxeKFgibv75v/TXqvgBE17/gNrGfDnmjMeuA+7eLGxep82keFV9s5GM/Dq/yK0uA3ANBwjaL1hvg
unOCFVSnPODIOn6Qmi7+wH8at/m+DmjiF0zZNPpFmNQSSMcd+3/Aty4wZQomC2PmYslQpZgp2XbM
6js0VCRl/MeAQzZPXTDDdMTWcWJeusXRf3syQfvO1/+mwH6E8Z3xl4NY+ARGwLF6yFogAYWeeiKk
+V3xIJ7kczfFanTS8ldLF390q0P2EzqnPD4zLn/CwB0UmRx+KEc+jqoZ0cj8mcZs6pPGJVM9W6ZQ
fuh2VZUFnMn22JqY1hZ8G4HjppaNZva9MzbHs1F3Xaf2xuG/R38CDoX5MISJaKn359wHOda8GekE
t182RF3HE6/Dqd2Y8f69yH6Gpz0ob5yj3eAxjre3c1k1TclNUA+yRRrvbqB7W+7093vVcEsI0fqa
Is2kevc36LeqiX6jVlJkDMD0ABTNvvNaZfGmlHhPvB/lvnwmrunNlLbK/qXS61hjSbuWsfczUonc
v3p/TFhUXSHVtK6Jaz166zoGACiAlanjd/e/tiS/t6yRht+S6IKmrAL+0Mjrh0nofvkeJVgFuHik
4Wti895YB2vewb34UkHiHZHFz1OI5gVnU69FgRljvL0d6poExCgI51GYesMFMD12bX0sPTUAMsws
/23jURDHIqUpETy1fzisrHUSZrdT9FLps/Puam5xnnwAuhN/HRIqsex/OEAIvLizUfgWv7c+VxmS
HQtt6P+3E16aAdxXzh5NKWWiKql9anbWLrEGou3OWfnEM6el7uQO/2Ey7tmQkxiK5HBF8wM0vvAy
IIr81/b2nY+TPFdr7v9HQucwMRZeyFFZ/RnN7ZFqBTs0ESH1TCYdlvY+Ftj4JTGedHss9c6YSFYT
yBRAPyIFlGBQweaV0vfT5Bp1v2p4kmizDluhU6sBwrOFwih1MBeALu57c2RiBXy8mqZJ0l4tCwIc
bxHB/8HEdPH8qDiup2IIaCv+s+/ht5iLE8+FlSCHPNaLLOlZLyRArwFEtZl0ZWQ0bmlGctkeyZBw
Tfvz3HvROiBUUPf6d7rRUX6Zd2aA52N2YQWGhIx0QHWQtVjKW3kzKQfn8ILBxfpCHuilrE11eHfk
T+zK1rTOrqsqQi6LmvWSA9Q0JkDrcTWdwTp/L+1LD02M8gUFrSV2oVueD70MsAgNMTWYxo62TwLH
HriPxqoPJDtW0Qn6BIAiPjyBk85awWkBbRhj71Bzb/cG8m/Y9y7AKPOJ9uwXq5j0KBqWE6TxKX22
v+CvThkcgpZk3wHkugGNC6Bz7AO73+nrSVjsRplDsQ4PlKTnf257m2kaFaC5qOPOxNdu69aICnFz
7jRF9vu45BTRPjcFOYzjw4ihOr1ncyj5JURq13jKmTJqUVXgp54yCZfHpS7kuft8MNehybfP4ngh
PC5Tsu7+3VKP5tatL4DkZizeZ5kH6Lz0QuigBdlGYcUAoKSc2PN7mS48ZG/CUH/fnvrAIr53XAJA
fZ9F1JUOXUbCe71ozQreBbLK1UIbSLtYL/SQYmmBhcFE7upi6QpudDHe9epR9LHddcy9EmqD1ZCw
ZuSLCrAy6fNuU0wyiw1u7HeJhDZYaMJQx+R9F++pEf4bP9pumaiJ+Ze0wJHEe2/A1eOcoxBDX4Ct
ErxeCtlyCMdCU4P+ghtAqhustaQU0v/Rlu0D1ddzh6O0GVgoJM1jtYGZ2trW1Di84A6W88LwhrIw
lCRjz/anAy8Wt+VymNpXadxbXhniikXQzfD/UHI3bVP3W37y1x9iKvvdodLZ2L/JGyV2JGXrw3Hk
8sshLNgxBmQf8y53uNjo/+Q5P+L1U5HYJPKBMzM42VzHxUQQaBze4m1388v3oLzKl3Kc4p+CsfUR
TI1ghUz5QPIhWHLalUtjap2Tj0dOeK5gTIbv3nvWycDXkNG4Cehoo7/IUTDxqe+AZhZP/E1e/UkA
ykO20qYMYLFVlzRWhAafdCXhvJ35DHteT5GzQVrA9d3gQwLjF087VKDvLHSmLHnto1q6ZY+dU342
0N2ILMnw7hM5p/3VKlqeaNRXBsXniUol7Efv3bAKcEymiF6Rt4J8yG6wqfE+0pOVWfPqVV8NS0w8
+8U9xhnLvV9pv6k9l8ghkdj882XeWtfjaU1cU8FDRqHAEODZ4REPYZxWM2etZSKtQLBC3rHan7J9
Ae96DSJW7iGht9kvC9XpBp/Q22soYVH1XYV0tTKQc0JLAlHRAyvsVepw5Fy9NI/MFKcyjalKt9h7
jzgjW62M2gBM9URMujrVeo5vAFInZLGEtgqPSQK1EWz6kAA6NrggHBIHsN7OuKw8Cmxkq8k4rHR6
c7D9tgycp93SBN1nLITQP8DOiH7RijTRXa9m6CJXV5XwZlDjiaXUpGGbpLFMUtzLkEa4QCqVhrpB
BMlOHCvD+agYW+mstKpLp/TeEBaynMNzFUwyUqmcAPOsL0ys8n0wqbj34nPa841eJXJFqLunIjk1
Fs0vVEhwyzeW8AEzyj8EtoX38gHHsLg+XmvWkylnSp8Tv0qrmldLhuEX19q3UnGUUDelF4ZWLxrW
NmQ7iYL0loY36lD2exb1TCvhd1/rAHEL6m0rZCywnQbAktrdnIIbreEcpJNiMqyH9kB/oKpKSggC
Ggiq3zAqvhGbX7PnU+H000fo76MEKecz2eKOQcxKetLNDDlQ/NvkMBkRJ246IN++Arfyh6uTdYHa
rpZMWuW2ptpOTaECdPESRDhSWU4Yd0z8h7WE08ex+7vwxb+V6Ts+vzK9V6ENkZTCaPsmV5v7Y9Vo
QWdu/KDKjbQ1rgI+cO7WMNuu/6mG3YPRssWHoF/F9zpVw9gWnfn0xUgsMnfNMpaPwNfZb/tyBLJG
AR8qjWUfjwV9BSF8Wpbt2mmXKExAQxH502QBBLjL17oPOiLkGJqgOPYUnCS6mJ2y96WBTrr91HEy
DfSyh67MnDKRayuTuuJ5RdH7B0c4t47iBL5LU7qtVc7y/JaozFIbRyCFqd4oEv8H7FAkq1k9KCjq
Tvnes2q36g5yM1fFsRmA5XQtRlvFF5SikMwdBJXOKZKhK7IuwZvWINnGgmp5Rxop9/IogcaftBpd
PAb1ByJBAQ2qfwBqnHDRsoT5O/U3nmFZ+AuMPOifK+G1EaBQsnmXUkauVDVn2MmT2+kzEXVDd8L1
pB1K43qUtI0tQkdPubHBiKxkO7Zl+nbJj7HeTiQlFoexBQxio7tQqvm7+YcMblN8LqzlesNbgpLq
ZlJfeqnX62Zf+eMXx5SSF6658OYNrSTPpWmATE5F2VMVJNIVkX17kqNXQLZOP/xAj+/tjLvBC5nX
vEp6yVVnrboGyZf/YZ/huBmM/bF5yibntJU6elxSwmCcDjzHXOy/t4ICYlwFXHwGSsOkxih+yRvR
OVuZdHY+/hPFDxY7/XSPK/TM2ABX8Rwi8lWcsJ00zNPvlFEnoLiCodgNlL0QYZF8pUqelTvxbweg
iZJTlO0aVRHrGxCGZ99I6FcWHV4AD0AGbAVaiJ+Y6enjZrfIq2x8tR6l57DVlYYFUuIZRpTipGj7
g48g46loSziLuI5T+P59/+XoXqDjwkKZVv+MCU5UDDT7TYwK3JONOI24WjX634ZF87y13O4TGjl7
x5u/pp7yPVLXNyOF6Na/hSbRxCjWoH0FbYAUKFwCaWHOA2u082Qiqsds1zP3kSoGLKChhNl1EKMm
uM+pVTKui0UPTxe5rQQUF2kRyQfnDF6Y0SkE06vigLUEeltYAoPgiCMNht3IfZ3U9TKHPO9teZVE
ci4KZtGHu2h61ZpzqHrGKcoAAUDda1WfyPawevvXmW1R129t5UCYFVWuze8l5cWywn5rG4yYEQ7f
EsUPSDQA0nLu9PR5UKvnQY7kmt8LapetT6gdUpa2HYVT3/Gao9o0P46PIDu/3zCPuNXGQMzwpVnN
EzI9MRoQ4VrKlj1uXLM71WdTclA7sVn1sZt/14fQFvXQV8fuItq19ECCzVm1ThmavOeQpbFsrJ1E
UlXV2lpHkkZ6hkralMmU5Q3irjraBQDFLG6BK8cM8KhF2Qkrwki2+3jhFOIz4kRBlaItxMplzh8O
pVpZLA6UWzcb2zMxIyw0/R5ZoaDlaZPkEziEgzSFgTqm9aGhpOZ6lJhoxRfR3e52iotHxJnXGmOp
s144BBY4Pox9o2HudMVY87/rIE4QlXiHC0z1IqQrjx2bLuOuyYrV4e4ZM1NnH8PJpBb5zOh2K2yl
8dH4wo4/8e6AGDNnUOp5AP2XHNN78r16UIfFlnZkDfJZdOWwJnjn2j4KSa0CsVyz75nujRas0XnH
GiiuwGFt4TaJ9McXi7XMIDfa386lonGoK+m6hJGKK7vMsKBjmP19hQI2TDpA9BxTHTEpToTGTNBJ
5HVe6kkJfRpK3YqmJiWPR1wmyemK0+s9jxNUmktbOnccqusktgTeBMgKaib9quNKbHbSVffbpLkT
UZjL8CwxEUKpFNAnrTmoFe1iDJPNXcNPtwuz+FpXOmm6vyoZltuLQ1T8fRxXqoynijowgGKvFdBN
LxTa70g3U2WtVxt44mxR5WkwFptnvrXA3L/+rwFMVX8G+LcZp7xtuCynzGM9oblIoNbptoqUPbdW
l4HNawXienZB7U8JMd4cizQql+F9b8/huS1+qVj/ml0neFDttkzZPTpgUiMArHegIkOK3V1klV6B
xHLWixX+oi4LfPDIG3NuIrmY8K0Y97Pjylv7UsuXmmohZc5wIS6qn6xR97vTOeaoLq7QeHmkP3aB
7oVhM8aI7hMRB3b3/ZE6PdY/YdrH7YBqYmtszrfp1z2SVuGvOr9T81MtnOU2sJVdan8M2y/Jmk2h
nU6Qu0ybtBhcWRjOom6npPUWZTz24iab/AdtO7qrqOIIA8wNflr6Ek5pfROjmS19oponDQX+XKk5
+lZpBSDTMGSPqmucUCezOgvVW3jH3YJOYDfuTSm+Ol/04cmwCBXjap80P2dgk2EeJc0zCuCPx0sj
B2wnhJ5VYa2VvBCVyMZSfuWhh9WAddqW2CNN24lKTj0JSHYkmk35YZZUkiBbvbcOg6lnXvhXSbLp
Tp1ORFUOjzylJ6sswj+qJYkhHgQ2DxAydazQyIKZybKWLB5Dp2cjDxiu92h4BvucxQN/TuwUri/x
u8u46Sot7amt6jwaK83mflQ5AbCoaCkM/lshDInQmzsMAhE+1e0h5/uZSQ3Rg0g5mjt+B8PXJhhY
mf8IcTsPj1pbtAUwjlAqSKIgMKOuXkG0DjAb2N2EcHUwOF+pa5MB1hh66slyez0xvBbwBhoIkMKi
/+i8zXo2eELFv2v4FFlHQubSXyy4K/tpBdVIiGpv/OFLkVb+SlUsL/X3wJM7FCQUZpHuSZVZetrR
fIFNimk9i1ivh/t6gM96DSWUJ6fHU1DM/3OSNjSOOTvO9ehPALJ92mtFsIq9oaBbQUCyVkJl2+ut
g2lRFfySriEZjaNt4YyU5BUH0pHVXclElkwrymnacwgbM+3XLKt9CDHpfbEVSmep06I8sFm9OhfP
fkGf1HR/f8Fq6tnlwE9QBES+UMIC4ZJHH88V6lcOaBAzwulzqPe3vgCVIisNqOHJntvA89AF5hvz
+QfqkYa0Zz1/fhW98IKiWbb9sP1f1/B5WTzEMTsbaftek+zWlRSdHjTYmui4kGrd82c4ggi40Vdc
86oMewyR0WjskegsxGerVCOl4+hiMurHiNlNoU1abQnXFNrscvUuGZfOFeGh+gSNE2yHKpXMGCEL
WiSXhuwr9ON5hCF1qnI36KKqbAlKY9Hrcjls4Vc3qkkKMlknBXoa+ggFs1uGjWzYXOA2q8HnqA/o
Bmo5UTJ0e+PINfp7szqyhvhPsNwO8foHjkv4UUMKcsn2aQNC3WAsLM8aShjpA9P/yhyVec/gGyHU
DBfas8IqASXdE5lfFqNb8BLdjPSzinbzwtCTeeQqM8sbNOJJNnqNKoqPDvKxunLpghMTZOcgguut
WuMZFcI0apOmwUhKIDJf6YbAXWGHW3Slh17SybFbtAlLZItPzRwAdAlNoeolTJVFSAWWbYbKDQcV
JDpf3YGWhRjY0r90VMsQLy6iURE/qn5BXficQj3cqKF59yc2OSl0zx1lPavSck96ObCJUHbCS/s0
mc/BS4k9Qey8Qju01K60nxEQBM2PnEXvSLIoz5f3Kkta12bfiuayWgVjzr46LreJzlu6ou1U/Iiy
LSN4kxpqM4rkjJxice7Whcrjm+lXT0s6qmSA/eAgPIbsDQSMCGZWUjlj+f/CuBjzJO0eckzvpXF8
W3B7sNlXKmmFR4g0v9ZeEj2+oiWYzXT+dQwruNzV8PbKzgSXc6qOSt4iM6OXenIfOuiet98SGnBM
LpfSO+OENdBwbicJO2j3w0ADRKL6d9kovl/XAXlWkM4MpE/2cCLpYYLfh5xgwgXPGiOtKZJOp+cw
NF3GNhKGabRYNS0ulHYZDudt1N5+OUZz8uy6kj5+gXwzpg6qsC+FRAF2aYX4aXqAF3ulqNSTNxBo
Fl+fdYZTTT5Tr6V88ROhrUuL9eBdLleDPIAuNOKedlNmg3gkqt55c+tAGC0JYDqsLPmvNjbM5C64
MjZtVJz6mkRuvwN/TjWcdaIN+/eObGEx4nTbcvRKsdei8DiZdHMgPhr9mt6JLzBzAZ/F2IyRbajw
URVpytvVSzBFk59Khbj7qRfYSOdCc3HsN1dKMH97aCRVOIl1NnDofW3pJUMZ5ZbU/uaT+Sv6fOgI
khR8HK6KqLfq7zdu/HTC4gHb1oSJVTSRTsFZmPVWbiYBcA4RjBhriDeNrTBLfYYFvh9zx5NEIFIK
L4THhF6T3eJLbO5G0OpceCLWNpzJkE81nDcSYLLiqlcRiXiE3kkU+c8/Jo146WU6oa2u1CrVd4HO
yQEG0l8JFqH+tg52HLZD4sBXFwKW9NTtv7dztFoROaGQBphZ87YOSuOwVy/xJ2eixP64B0fUf5qo
jcrwsermY4ics/961Qzd6qaE75eWRt1nRN3oILzXurjP9ouyqWDp3iybJQcwcg4Znc4gHl2/GWej
xKlcMyrTL7cw8CqelWlFDPYJBlKGqBUdWY2ym9gcjKIZEgjpj+Ae98FYRYpa2gRJoheufR0Xcs8W
bMjsvB0mVTsv1fufoQJOPedR18mZnF3op3JLOn3AkEV/3y6bDBEYnP7ZULjLCA1tvO0Zilg6V/Z/
QoFhxBsW7DQtZty90ClWe+n0Rck/bU9uzUWIMrEBPMwTYcDqFRih9XtY/GiZxJib/0I1UkOSargL
nYrKEj37uGsj/AfFIE3ZGsKpH7iIbWQmg1aUBe2f/tNkgJZT3W9jaUrU6UAJobBgWkbX9wodC+2K
SZeuiGPDckaEwEN86jdEGgJIK1T6A4pgYl1G14UiV/sfB5IXtybyfvMiZ1Nd0g+iLGb63qUNgzYe
CSs796SVIsju5gPfGS745T2HwmkPoLkUIaH68NOzc4bOpEs+39x+X+1ncmm96S4jeACBzJduqUaI
cwdYD/aLzBhFIq76ZDcehwbc0c0Yr3QYr5uXKenhtNxxVGTWSJQ1Rgsi2WVQm/OYZ0kS82qtf5rP
ETs1Ok6wnKkXJCrdLYP+rOb5r1pHUspW9/G1yK0p4AZKlkBq2VJnDEA7eQbMtKi/PaTmhv9Juvxo
rRGSsi53qp6ELnr3X9LEY+mr2BkU07Pbtyv0ad8rcI6L3cP0ibQn0Yi8AgNAQ3FKjTolZXJ9erCt
/pN45LLZqNa+qVYdXO/h2aj0Cfo/Ib5g9L5G4MHNsrwmC6aBJw0O4DGBNLq1EBB26tG6udKzNMhF
Qx1pTzl4xvN/PlnXN4Zs6dNYjKR8koEJs0d26dHUnVf7J+BgqwnRU0h32sCkIsxUCT/OQ1kJN/f8
91j4uWKgHe1bwBW9K28EnkPizF43Zm2Gr9baq3gC2owFFadYhmJ0g2W2CwoegKV2d4B+1B4A3GnE
ghYEokwp95GckH0kJoahq93rH51kG+Bm23ngocbsEVYR1mkA2neGj8YP2YVEKbZzmp12+2+boxIs
HaNSm6zBpGLux8RVp1823ro1xA24eZm5HYvOt9gN1R1ZdxHesuHuXGirnBTQzj04nZoT8V3Nn52+
TrByPZJat3jwWsnma8nHHb64PB6p/wwdnA4zdxafkX0GRWQkCdxi1k0Fla7vseYHouogko8veJB/
LGX2uoNwogH2W8ynYsjl0MTvnHxKYe42gcUrATICWTcBIrqIZsr8OVoLssuCVEdY2DQREkGACD3M
pOgWkFHycsDiyq45l433CLZtuFI+0CU4I092tgKsatqJjHFTxl76Ic5Ncp/VenZLuWq5s4NED+vO
zHJaYUPhJdLk+7sKF3wsTqu8HNuPDYUw1Sw0cCKDBjevQNdcBypcklt0KvGQd3auqlkNQufRd7Z1
+LwvvD0WlDhrmBMNk79smQmGYXqK8zzNhrGu09YaI3qfzaZVQtWnLM/BlYLlMCYbxhUwbWpJ8gzn
pGH7Pdgp4GRwKJz1GxV2JKabEfbpcXF+VlBybzqkrncz57VnjhkqgdFi82Z9iXrWYpKOfTBze0HB
9lrxJ1Z4SU6eKcLB5RsqLBM5TneynsiLRHlW1sfsl2g15qSGvUkC/LZ2uaDRQ7z9AE+0DmyHwMIB
RXPx8pulBOe3WNu9OT972bYfXl8SgBAB5239znhK8Boa3n0d4PWMhS0yPIWi9jNNDUU8Z0jftdtA
2DCaIJlAYLaKrEEq/gK8ODFVY0MOucJhW9dl2egG4S5oO8S+Mi8X37iFbO9Hrk+e7UgiQIJQ5eSg
MHhzQXFgNtOXvCv2nIfzs6WGvGFCF/kz3uR+7dXJGX2bp6hXqtJZy9TVlrD8hpvsWKEnAZFvGLaU
lhaFYHktfpzd4o6UpgLVdAvqRZpbDoW1MkLTjJCv+BIyJTVuo/vie2mvP/Evqd9rXP0+mkOPVH/9
KExS5ep8jRT/6sjq78RK/2+8xWd1JVRTzG6HQ3XON58sd4vi6gOWLOfoU6Nj0aW7t4tXGQg3/3MB
yK1j9Gbg9zZXxD0Vm3d5CZni3x68aSBtS7oIxsP6ij4/aEjv14N5Z6KKrBwFAadV9V8rJhB0O6Vw
zsUc0IkHOV8BrBKzwyVd1Dkk+14LZoAufFi9McLRzXNRwdxXzDc+/k7Vk9GQGEtw/yvbeuWAFkys
kt/IdgcysETkciiTilxggwqa93XjyDW0GGhqRiOux+nQta5z59gJso3BSpJIRdY1DLdWrLW+LMJv
MxjNzVdoz5VrK5+3QLMH12+P4W2W3ouLL8hWFcTjd1i++LoNlqV01INbGxekxasYfggIJOaa4jUI
7Xi4Ox0RpvTK+pep2MwZgcWidSPVkaMIIillKm78/xqEKvMVwDjmazGniBoAlQ5UX5jighF4NfoN
EAlCqzxobZZzXgDyoCLOCDeoSNQg4ZKLGppCsw7JGy7gXCOLxQzTMIQXyd84ziBAEIbd1z/2/apL
SWyOrYqNFnvQnyPz96j8ys5XeMBYaWE6JJWJGANkgEOQffoPGzTfj2sbn3TiXmAtpL9WXC39dTiN
lkXse4D3MT8dYmNAmcW8InhsL6k/yKGU5wexLoLACtEXCzG/+Qgm2h+JOjhXa9qGgC2xScUr/QO2
waSysrqgxWBJBW/d34Pu1jioZEcxLW2tpmPTe0K8sViGIOHMFP7IRH2eLsXsqSX8BP5NaFNGzVdR
MmFtILUADISiifq/4ef0pV2vvSBN1R1FGpAygeeYf94xeG5mDucJw0O2zWNSWtBMxluMcHVz785J
lL4juklJLddyF7o2PmXaC0Ve0up9NbVcj8uR66ktZSJoShn4AvzvvkGWLWBWExc31SphyewwprGj
yUTApaoui9tIBBYvQ1nJP481SIzDTZC2HB5AW69gmWLgkdhj28NJqVPZoHtBerIivNRpQ5YQgam1
rQ9ft1IzCupbsfsA9LHq1005HLE7sPuJBqxW9CaRV/+IytgqhgbMwxY8duUpKUBHAK5Hhy33oj71
B/DH6MW4Rbuc43d9QAfdEZ7/cqvxPQDXk0lI8r34QHtIpcHWik8XU47OXR2OLCqFyW5dmg+YtiNd
PyWoBIqcznnYnYE2CeJiz+XphlisU+4w0XmBNDHs5kO0ybbnD+jBI7LK7XYZZkIOCvRbOOj6nEZO
80EmyyIZeNHz5PG5+l4UPRHiXYJtmfmq9ImkDcp6ztszPZYBAIYor7f9MjOdZuIdSSLhQwEbBzcs
JiQl4ricxuFLzxHSNtXv2Q/vkQMYJ7vE18jJE2Og7PLbzZ8v2Ykq7SCDlb9Qp4cOCJ4RUqfEjS14
lYl6ELb8dvGFbBbupF27oLXSI4cHH9S4JL5qbRRM/yCdF5uT1yr5mv68Shp/YcapbAUi0GXHqUkO
vhdd6KiCjNVcdUOlYsQqMSaf9mpTNHaOWbY8aAFdXNIJqWXUWdwFADh/MlP5uxCWxoZD+nQrC4Me
SlJn2pePJFRO6tNSHkpm4jnDym+PH9Bv73iQXO7u/R/0lmHOWEVyNf1fIYncnhexqK0QtkV2yPPF
H/IrtlnmfhRuZONFdGk3iVKKclBBwZJixtuWOFIv1wE9DpWgUVwTdkTu51As9FzH6WzrLmk6kFzB
1zBOv+7DZ3bGRS00jeAYqYfKzTQd8rQnsHT0Fz5KKQf3MjdL61WYyQmvJrfJqJOmaYiueJQ/cMew
O/ddavdWyNfY+0CeoJQydc+cZERBE+Mc28+sB+TR888m+wS0XL9UvhTmyNygyd166vFzeIigTvDI
+UZoL/2tNimq5sxS3b0zebuiWSjLT9qoFCjZ5Ac/a1hCMqQ7vPHEw3fCSsf4Nrg5GBZDe8TLbvHy
ui/hMV6PQF4JrXt/NeryaHBSCl177AecLEp0Tr8igshKcB9JoOIifqOY8BiTkzkHEJVACjxK3ht2
b+IoYKWBsYfc/WsCuZZocEE23TP1fYoBHQXW0Lwn84QXFqXn73wI9vaOAHkEn/9CgzgSglJo2drs
cEbb1Gxb88DKWKUn/+6U8FoV7u6JDQpa107/YxTPze37hDQMy3fBhC3rsYA9ht1D/OiJekIHRgzF
n05R4lmTVE6fNVRiGqMma2HtL6BTsUgw1/8IIUYLRa9v53wzgq+hq9grSfxt4ZKaAkWR5MGH8V2M
n8p9hQbGgklcVUYuVA5EUB7SXrgiaslNiunYgvYfV4pYswqv3MZpBhGzGdsIpDwhky3ei73mve6G
dQpggAGshqAuKmUGAI5XF5bhFSOS6Eat4TXj5yXLMNs5PvtB76nMsGRKSkjQF7+X9lGWKuwJmTDU
/tSyBRdXpp+0VszQG300yBHgI6CvzlzWQcHfbdRiATnGBk9UA7O+la57xoDwBVqSyzfZWhK4zivK
HujXmqwbpbqIXyh5A4dE2xHGnLxZsxHK+9CyyVhVjINLUgPyj2Or8x908WZkoq6yd5IIplY7X5Y4
CcOUKCExCtssjIZTbm+798vfOpJYpyZa7EAPFlaUH1CHqudSfYBrAo34fCFu2O9NHf987C5EFZbQ
IdYcODG7B2JTfluYRlVaBsl3Xer1G/f1O2f8+GbNc0m5rfTWzGhJeCv7F+nVi22d6esC4W53qM1N
hV98ZXK0TGxuJRU1agrsurbmdrPhcMPq6FLbFVAnDRG2LfNSY9Ljmx2wuw3fzn2QcTORiH5uu1MC
Fk7mZZl9YegNc1S6CIrwxzJ8vPra8DgGbdW5xXU42dsUkaf8Odzkm3tp5aNjn/3LKJFtnJhciIpX
ZjDEFHRQiPm2m8F1eZL5xdaktWz+ZELTip+SGbyHaf0Oyx5q5uQo40QN8MUqHBqw59nXKxjmLhx6
fJbPBk9QtqvL8vbOUH80wkhtf6jsbMk9meOUmlbsXdnqYHXSXwfz+aScrxKGdYHT4B6+O/jhXXZV
k7UIFgrSHUM6g5I2i8DkKNly85cGzpU7TMR2FzvvVX6nVQd9QMPnz+trPMvufjOrF8zHwliraVii
4P+fChXZNBviiwUp6pmI65ccCAho3pA/yYHv1YVSbfb5np+v8K2Vw40b4ddvwwmvfsWJpVn7SeP0
hM/05AjJ7iHB9ojbA80rxdZI/+qRBZPCcY2XQwi48FPS16GyUUj9+/cmNpjtPUVjBYGhozH0b0Py
0jmiQPx5VSVrv+WudEk5kW9WtC1o9mg9Ywilt20jQEOUM5t+ic9fTPHX/1X3NUdaHEvJFh8HjYIT
mnLbfzGlU8a82/pv8+oJYu0dkXVZGX15NoiQlta+soogARxIctXYQe5ycu3SoRYCoHxs1IqZoiv7
JN/4wlEro23kgLF9by7LdWz/0jjjdnlm2pydUeeMMxuWAcifZTwdKjXgZ8JuiybE8gBXaaXiqYZp
4ctTxu2tpAmF4kUnHGavWln0ThPirMbb7vttQbekrpTGRBoQik4KJyt44rC9q4tysVxvTJpb2kn1
SH8Vifs/s639oPlBPWjiKPwIlOuGSQIV/FO30B68CB5dhg/J3mCYPB1Mhy0rYvr+XkHJZ3buSYLq
W7F47eZVelZw81sFcSLtLie8bvLSnqS2sUpBJj/Z76Vr92UDQL+IJZaHJkrt48wALfwuehPTb+pq
kRs60taKKK4Dc2LmhQR5hUvl4xWisUY5+S1a4RLt0vJ5cl1Bkl0+tcO9Gud83qRnwx5hmxcEEipW
VP1/inBVwdo2oEgEMSdoMCodslstrB36iMj1TgLfu7dKI6+AZxgSMq67plhk+LgLMRGr7vW0SFHW
D/D0l59Gh3557dLnrKa/Gc+oWjLoOxvL9XKj7dN7x94t5YLgvOJdsr1bxXjmbXzlHXShLLEYb68j
IhK9JPdoxu80oc1KjnxE5PZVCENqJjvcuZmhAGD3eHWDNZCsIIpV5IFMgVIt+kJ8Vc6iyKUnVq96
EINfZMxcBk0+Ay3aMUEbZsWFIcH2xqHvhrXNs8yk0FpBg35pb2JFTY1iP1mHwIvQpznKcRNTIEtf
ZJGeyz70VqVWvl7lN0VWQQPdmLqeLVwbKSWMARvnC1QE5EdlPbWIti4EU8mSI8eYvUQYz2vWRq6F
brWRe0BEkPwrwfkyMKMNyyuQQ77O7UqjWhz8GdzOu52AiA7LIRFeXr9y+hf/0on2jRIu/PXBworm
zXM/pS41XTEb3ETDxwHMfiBgtyQ7zbl8zLN7+ZqF6xxD+sW59OCF9CC/s2j9sP6Cvem7FChMIU2K
TmEKHF4jrqZ7qlM7WZ9FoerhPrDfOnIlm+9reDftAw+hL+3Ma9rtJg5uIiKCBaL/7Z4B4tkx52wp
F1sA0E8XYpDbwW2uvI/v44fq0HPN4PiY5fSe7QIcyp2SOSD/J4A9xPkintdSH0ltPO0i9I/eDa8d
NzZ65eSFwbD2iHr37Z25RfoJTA891B4b4Pkbl4geuJqvFq5fYnW0q0R0t3eTgxMnegeH8nCpKlls
6aLgSJzr40MKCqa2TWx7qeGWRzeUHsMzf0OPrD/OQ0oNr22ELOwQbjn7mSPLNW+L01mpW0e4hTJr
/AANpkHprGSOKNRwPwplWO3Z5N3KPDn+KNEvsCo+0Oo3w+kPzarN2nV+iq1RE0GJriSS4bjK6/fX
noEsJx76oflJ7TNYISzX5v3WAU39PpRWVuJhR0cygMrVKa6cujcOwMJ+uBq5GVFnASCRScnSasK/
r2rM5EBQ/8rc5no/dC5/r9oLPrZX40tTLhrXpMifGaUS2mpgh/jY8mryC41hREs+yCg0m0t3Ljsq
3NmScs4vlGhBDCiRzHx1cGWYkCvqTce4nw3nBd6THmXSshLclmjO5rByRUS2K+OC7AhjFLmhF2qv
3SLjByiOnZVLmLmC6/drOvz9bXauVsEghtMrMRP5eT0rna5YemPQ2Kx+pX2ZBc3O/Gy+pKET8Evc
ieA0AOZWoIuXxHz56IAoJDm88GTSMp0zmzIOmyqOJ8crwCfhZh9awvp3Snt4OU6dEAI//YKm7z8N
/2VKSSGuZ9AKyGRRK04FZGlJxxjHFK6WM6Yef1VQQvLFOUkKUfjqLwpH4RDAhb0715/ynQxmKgVo
nn0cvu31ylc+t3jbGZALIufbrHQmKJ2Fqk/f5qn4rZNwvhB7gwg9hz2n+APZtSU3kFpSgVwpK8v4
YCG1BQ7YNi61Xrk7YQSFqVft/91gxyD5j5pEAjQa585wRErrjpDxsLmDOkms+5evN+vCG3OiRcet
GsFY2zR4JtIi7gbhy1vxsqk3rgTUuWIyyCDsQ0Tye3oLGG3M48oX5zoKb4we05sF31FoPsfQLZiw
jB3iq57P4ln741JNr5fWuwTsBL11UFIPjQiWqF816toYuNG9dn1A7+mwYbNXQPwUIt9owTt4JtFI
56qcy8t1QwnrqTim5QL5RdnmLzy1TykSN/R/dFc5v3oDaiqKZumKY0wrxnGVJ9oL9+aClDUXS1yw
J9cKUL63PjX+I+K5tOwa/JALAfmD/ayO6BjNhMdaPQYQuwUlWiPiyFzNftY/qYgBSSuspLJHyrm9
91Ig4k8sKGjIO0kVnRGcVM8LbJj2jiUhroqpyoAfyrXNuZdosZrCWZf6MItvUSCTa6YrjERkQJMn
lguVPkjcvLrFj63H0ifsG8XXxU6Fl9gUHSTxewQIaKA52zQd7C295+OzbAnt6D5ayWjYgVES14rX
oKYQLFoJ5R3j7T8+22jss2oE9J/HL3CfQiURuo3H1oicXciG1AT1QThRwDDaQJxM0W3fzjGFggMe
Nv82U8DN2/jXqXkGlCyrsc/wnyFQM41zq/1km7PfCcF9Xm6xNGap2c9pSONUorCev78q2HDI+/cg
CGtH2UtDsD3Y/ETE/FP/AMqFOGX5VRdtNxMfu+iMMJF/FQ9z1FnukSP+jnKijiQMbNCi9DNMun5z
N6b6uzA/m6pp8R5aXASdV2zIP80DDjpHIrGkZzoypVoXpTApiCH1AXwfthi75fox4QSdpV2YysdU
uIKIPbJzXUWZgy9/k9R4j0TZZ87MAIp4TmTbXGuvi0f5KKxbN25LmO0MN0QcoennzcV3mmkvXp/v
Ic+AIldiBHlp2DWU/55v/0JIFozyr8zT+4tLm5e8RDoocJAcKfYvTJQyyENymcIEgZVcAcqakkpZ
iunG69kpF8qGt5oxHpkHTMOOB33Ft0rcDY//OSjZjIUB+1Jc97zsefiZ+K9DgcDXovmt1ENIpVe7
aP04G9hWRtMJrzXX7fX/fA0ZfLOgQEz8n7LLn7HVT1EsJOXm5TszGnuGrOtOuJ1nmI3dQisJKK+G
AmMgpfqT5Hl7VvdFpJYy7KzCZ5lMXCu89RZyljUPrPj2gQjPvm9YKLPOJh4STYwEWh9/SZJQd7Tp
YjZVXeHP0t+46VTEP1T22hMwfR4DRXYWWlzugGVqeoAsF2kM2ANg9vuzhuulw8KCO5FiaQv+qFSN
iavSeCkSal7iWKfRpXoI+xqKOXa88e/l0n88xQILWO4KjxFpYsuDPLFJwCfukZRg53uRK6QN5Bf9
AjVbr4dQDgjgPnzGvP4WSNt95nCvfv0B4TEbO1AjzmTUE80Pi4PJIktA//qeIGkw6+q8ch0tPiLF
zjw+xvQSlnQuJgUp1Akuh5u0sHnHpQTpvrgzJ64PrWvyxmvSL6w2eq1m7gC5KIsR/XAaGC/1t88n
YUqd+OUYOirSiG7noGXjtfxfcVLXLD6Hcb1pnQtFeGauhNB8lsl35pUAjoWSXsom4LoKfvX1kA/p
HFy6ZWeRClzQ8l70RwB9l2WgophMb7kKE9Bzwv9GFgYb6a02kBw15FmnDmbCLW3GCYvLkQhXwWX4
CnGckPy7oyUG5Ivxc6JN7+EF4QeoJzcAF9mrfLV63942nXRNUz0Y7h1kJLAS+RWghnAJ5imMJ4c1
3pJKtCdGxwOHdLiBzy2ZClMxVCqhTXGjv2x79gLuOHz17d69UI8NwzYP2CKfL45v05+QLXuo7oZB
9aVIrqyR0g/KpqWVmSD9ElzwemxILFlFDfqq5RdgMRGHFJJzTBZFSQwfE+R7WIXPm+jgWCpF4NjL
an7T1o4PyTTMERkvoSH6J4bkpc582HSKD206sY6qUdcxWsmGC7fQBKxNnvr6QoxFxiTs9Zj7ZePP
WyoF6K/dGTfWR8+t0bvjlW2+7E8pudT8YsYIx5dEsGb6U0KvAX5P4M2C3Mz8EB3XZThPF5AVTHLP
L75NFqPZtXK1JDwdUN65+G+wkfUAYamah6OfDts1L5QSsnNaviPRZo/pGBZh+LZ5VJ6B/6ErAa0j
WWmUbTntttZlCT2FfWQcQNcgni2Y/N6e2ChsMrczDaP4nQxSjr0i+bwiw8exdeCthIjh4orJN8QL
rClqUvY+ub5OmGdg6Oeic67Okbppwi9HhUBw6bA/em1tvhmnyM5s5qaaBX3wvJG+ygJFxDfpu4EX
VztQs5Ol9696VTA+tsA4NSsOvzSi70YQPvgHmaRQTGLKq/72o1xPjYzXu5c4N4pNJ2qTCIvg4L37
fnLf1kYE5ERZUpivt9HaElSEMC9Pvru2FqkmDi7E7+jxUZeF4JlRlPVu72m95nSRPgvW/AQpHfNz
+/tNbRfVXXqbC39j+teficSwZ6Hqspl/KjcLsOa7gNzAU1uHHNcEJlomEpeTMVL+j8iBeVmnS7Pn
F9PCyO/LcUO0Yh7LrDZv0w34Y9z0UyA+UI2h8lEQytIF5kSOAXqzPprqRTAvr1Cvq0Re7Q2B827p
L8wpGhSGMCP1sAaAaSGJ9lOZv/pVeBV5vrBmcL5HvU0Mmn5Tj3K335r7YD355RKHa9JdbamvveW2
CcjxmkFyvVN28xJCEmUP3YebBKRC8zdsdnGF51RPZvYpqczJe2bECZAjxeCMD5y599D9pnYOyaWb
wIHZ2twU9GYtLWVIGRu5m5AfCI7XEVOR/uE2prKiSU3NWvOAgxwLEoU/NjPEUpPDDLPV04PSVP2p
v6teRVy8NgtrXQZJEo+MEqCwcFTMIoXY7LgoPIPUBiHG4JApRZJBH8p64vA1GS7zc1aDkzbqk6x0
nQ7bYY1D1SZtHYz2efvkanhoG0fSeyYHIMOBRzqUpl1y+vn+jSJ5DHO75J97sIIsfGufxOLdfet0
+hffMZt2iNYPazZpD83GF/Bi7ihfw+F7zGX701pgw8cjM9ytAVPuD67ytp7l5rdT/O3o9qmHAyay
JXbtgrogsDpn9VV8TzVmHUVIEqElA4KH6f9aVwsuUPto8Y8g4c/emVcOfV6C7DEXVus4w0Oz2ou9
/1Ih6A34YiRQLryDpr389S9FGJKfH7bIBEQ+iU/RLyXeBmB6DUs3C9bhx7kj0DCsABs3tHnVlYkm
BP99TVmJODYb51GsVWYRfbsYQSHNDxWmzb7pEvbUMCYPJPemZiewbCEeoiNJ5cLZREbrhz2rc8PR
1YCzs2x8p1jX3rX9JjUQEACY5F4L8QZW8Q+d5E/U1gOh3nrKyho5EwJYoDNSV4jgfE2l/qxyuVO/
Eusl/3Du3w3GDH9UvwwzqiLTnXpqkH7odaRr2ye2XU9yWYz2F3WQV155RpaDOyuLmWrFjUdBJ7f9
y/CpMlsN/yBcHDoAvWr6CO8vuhldzoSvYtBtcpPTTtE/uSqw839s/GohzyqVJQGnau4yYtMRInby
qgZnx7uXowJ8pYpic5qef6b+b5NIA04Xl5qRpaGbLZ9BNHjfJ4ogpNuh6HOFWBb7y9jDn2aYjOo4
MwNyBeKi0a9QQLjMpwsnE4XKD9+PI66fLr/wt50KlvQJ6w2nw8axc+oui/lws8E+aiCKPF7sMQTn
kHsbqKvCVXazB4izeOKA6IawKqR+lStTLAbTvF1qT5R34s9zDW5p9M8Qi5yhovbCY8uoJwfYgfeq
aDqBK0DqjiBB/770SOK/DbJ/Ch+m/CDRWgtZGsvw1x9+tSn5GuUVY6YAR0vFLIsGK69kb9zEsk+F
st+LRdXPPt/zgDL6OyjgGFUmKiyNaZpXUkz3DzXE1jnSK5u3IS7J2sdKcnkR/jWVNe80AHqBY5cn
7HdiLmp8XNorV03WsVCHDhzaO8GNt5OSPhavmxm2n+daR2kN6yjTsQdyFFt90SvwgzkuTocUzelQ
XQq2vRvzYdIgWS3h7vQyuMOQrrjo3iJaFst2EPBzibVow253KA4SgnpYQTt59eFgRchPbirU+z8u
PzU0wRjbZorHzKKTz7Y6bJMG+1vwzyg7j9Xgd4jtHXftdRGkCtpSlDWUuuwQAOFIznILelAuIxkX
jFgjDK+cCVs9WtQDTWzi+FsD4vkwubg8bHG9+N75LyaSyCeSMg7s62CwrCvhgGsXIP4qDECJ9Vdo
kBUAzJVV1HfghSpL5Vm14im4obsLIE9aXYQVBRSma9pYF07ZbMpTlLPmnLVwczJ5GXbl1LjoU1YI
icISExGw+tXm6+kefiY6lhw7XiVV0tM4mAnJf0S7ZvlkDbW8mpcRwQeSuQ079+8+AP6YcjoETd8/
smyggdFmEawJ82YU/kQok9ufl2atX7NRXZRUljicIdHIfg1FIM0jM9cGZUrvrLqW69caYL1tgRw6
NfOZNui1DP66lCcDZMDCv/5BcqGRYvaa+tQ3+nUBgdzrPEc+WDMLsL2PhHCRtdB/3JiiGvH1vVSC
c1pOszCDmB8YiQSdiCRjBi5ZiyQiiR2ujPme98PLWM/6nMHwgNnEOY6edJ7PzhxWAobSiTOrosji
d5ZqGnIGylvykRRz8OW7isV7N2bCk/jkCp7czFHAvMZiUh+G5SHP2xIHiWGWtKaDkY1f2PDy1KFT
X0T4ekbwN72rTjlc8Y7C4klZ6YxPUyHrtjg80t10PIcLOPU6kMrTsiNMhnBaluIBKhxK21Kgq3pw
/7sXZoTJHhipuhHohpN+pGUnlJUeZFxTd49kgTSG7ppN2nQwroNVIOSIuL4EYdEHvwOmgCxmNM9E
tH84Ksi0KN94ulue0pJlguRC6y29bqAOlzofxqxi5t2OSsTs/oL/0LZ0fPyGPGGjQmCgTu7dibnj
UfDKno3XL+gNR8hUCeXaA45xW1X8pv+3r8ymwucOp3UrlITR+RuPKlq2frwPjgBSngJXwm943Fx7
r91zXlXdkOaLEHVpYJxaCR1QX/AgZdCfDNM4IEczTPpj9NZ78elICwmxK32ptna3DNzeRrNOUbza
nu6J+l+QHHozq7TqDE26zep8eu+Tl6StVGk2u8Oun4YGZgzbS1U2diuYyoOVhpYSNqM/bFMx+bP6
dZvAEGMTRYyd22YznDtxT1CviHUBuICu4O5eX22G1HalVuuyTstWCSWyel0aoFez0a/9Bum3UaZs
dhzDHeHtI1BBVfksd7gD0h1J8Nu8+jgV55gHs9CPu3K18813LNlP9UxFYwR1R/5lDOBw5sfJMPBp
4HZHD2er/o678oZZ0MSY2vs+skbrYGxV8fFZ4xZLZidoVzPrBJ0ALFH98fs+5U0qGnR4xpKB8XJk
2lgDSC1tASfb4aetS+YDARFes4m2g43rwpI8md3gaFMlBs1joNn3lKUoBo9NNG7QDtvdBMzezWTi
a1LtXqG8mdmqc5E/wYH0Q/M2n5q4lHd5EX95j0cCEP/upoclMGQ+ixir0u8hU/5ZqFaPQwncO18T
J1HmmDIQxaL+EhnINRLdK6WNMvgvIog+SVzKGlXubrJqLQwFthFYs9eLIrO/tdaRH3XwWA6mjmj4
/XQb2KoibU5xXY7CiVx06BYsxcMRH8UDn1YqDW5w2tdBfOPmYUh6w7FmTTtIAdLxBy6B8LCek/ZK
LAUk/SNM7V4Zg1pGnTOXGYr1oZ0qDaarSlZ9jBtBlm98BjR0DIo2nPS163bdeHhqgARgLRK7J8it
MN8lzzHNLPSQT3TeELflfEf6CHBcJc1iLaPSmng1RIYq5mGnLhxqzaLgEXZ/sFbDhAduT5CFRcDs
j7Y+zSK9LLrXaO98HBT6QpE0Xciw1UCPQuc5drc0FBGR7bSuQqHwiCoprmgUr4aLdO4iuxN8jQgz
tbKubO2B0W97NUqWhb1IKx/c3slod/1/XF3jmsMYrPboyhFzM87XP7Jx4Ry/IzzzbegXWYkwwv7C
Bf882lwpgXDhPTvIEse4I1pu3xhrpiVpv1EpBw/mDhyXjPKtwl3YX+dy6bm5R3x5MFc6bj/v49Ig
SeVE2ldpmXIyUpfpVyA+LxI/AecPZ7PcObGLj6d6s+ym8sdgDvRMnc4SS0xW0reZ3idct3v/HfBa
qCPIfpnBfcEtWeAwVm0OdobxW97Crzl2vMnkjJIgnXPy8qsoSJJ2a22RcEbOLARdZTOJmt48hC4y
gkei865FQfokb2FTb3S8BYrs32mYg6FwX8WKRqOEFpWnNLtWR33/JiqcTfj61SrxtfM8tkQdQjpW
18l36+vS2zdKVako28ypTXrnvC6KIPO0r8RqdgHvpxQyJYnzRhpaO8YkkUYS9coWr2pAuSzKpxbB
C+NPHTui8BbtLeYP3FaIn5jUzb9xGG4kOchzqRXqUQHlW+clrB86Js0gGoJPJj2Lf/PlLLTxj0jb
KQBx/2kWLZnjff36CqW7OEv+fIGB0WxqadosPInXONmwku4bzx6PXAtGgxc7MM2k18tr1XfAtXae
OBPNcaGgUp9OnarjuABPvefSVOj2zWTFz++fy8Z5y38XHoRUVK7JD/wXanrbiWEC6PLozTFiHbhS
d1fozJIbV+BeTjH/+WTrtf9P/Fd3wP8fFkgWwjtn9W+HulIMUBUebneq9JG/v4IFHVfmOUFjJok8
Uyu/N/jNo6aBqPI/g+DervLGDKtiATiuq+APHo4TTF5wmLxbi4pUW0eDHVWZ+1qeahcgP2Tq1aDh
aXfoFZcW1hDtKgOjrM6ejsKL4TTVRaa82/TyCNA16WrtKprGy4JCQ7AWD95npuOhdFBQpGVLN4sh
PwEqVLNVLcz8KIv8y9K5dYnCwUarXNcxJx/zNfOTS+w0pkEltvurqFwTvG7EAbGAj+s8gJ1BG68A
vB57K+loYen7DW5nFi+KjIlmvbMHGAGSLvkZdSGydo9nuk5goeSuhCEABa3gmREkGkMm8Ggcw6FT
Dr09yCXzYDywhjkoVRp7W8aSiJZkyoAvx/7yEKCV52DDXgCytIGscEKiqUtqlqIcKgibrHDoCl6f
cyndAaxlzbweKuKuNGT7EUoaksZrEa1jm4zgk1iND+gyBMs8a16XaEuWVl2NkrpTil+Za+j+CP4J
U88dU/cJ9EfJlPTceuIAirJK7IDlQQCMGnwVZMM9b5jSuvBrs6fJ3jY78SQLbbNv03FEnugHPDz3
lmkrGN+aDmu0izzfirL1Stbk3In2CQMQUuzAZlMvFqfpbng7OpmtAqCDie5xmEkq4eznszUvGN/c
dQ0gTn1kmO5XCgfSakMwroHXiSkb9/yjffE7edbRjytLw/ONRF4VUMwjpEGA3VoQFcgaWu+0CkZF
4eV1TQqrC2dNAnUCntnEoDQz7GmfB3JSVoQOZ2Zdkm/33KMf61ffweRi4QHSOohy/6IeweJZqOJN
90b93ifUR4cJSsuzNj6UqjOUJdjD2Y1dmuS7QqBaQgjK16xSIWRJmCZd8Dl8kR23hZgg0wPgudKr
iucdrOeNBcl5HwRh9MVYHuI06PPh1nU0ohWm4c0jWcqI164sziVYVHK3JKsYC8PWaLCZvpsq4X4m
/tG2iivM171+otABEOA0dxuVKlyQx7sTcMyW7F1Ulg73SzOi+Ry1CLA3QwjSO1PzOgOQLpBU23kQ
BJsMFK4OyinRNkILKmFqByoRET9xGG4ARLo/jb7462IdMSA8PFOcj7mmY+d5WtZwF6HcdeqBMRWI
3qJ8H0eZVpYnhTmTs5JdEB6nrlbW96pmoU+9Puhct+/+eGhYB/fxuArL2oZ8s/9G1uNtTvZTvip+
6krss+OUopo6P/cxoAGZbNcGC/FWifM4IrMorkcUSMx/DExc5dr3H2NgeHEuDZgaCHJqC1BfY8fb
Mnf4rb9lSu0VMqezncwL92Z8a5vkwBC3qs08qJ/MuUBeWip13EqkjNX6zZ/8UthNAfmIqKRmE8Mz
oOX6RuRyTPahd5lT5V0KdAZjzXP3zVYXWcR9ExtVi+3ZMvv4stvyCvy1aCZg0aqwMBiQBnH8OEQQ
87Yip5d7mXRbIcSmmkWdYxvUCEvJbLoVLDnTUkATmj/wvzujBKuxhoVdxiombU1VrFRBj92Dm67K
ffDsIqPFlYRNULOAWOccF/57V83e7aV+E17MqxwVUNuu/ztzxBAIhKe1EH8DtW8DXMPQDKmAYICB
iWkSDzhDDopdk3uIf7Yb8Ml/wWmp5stG3ZyNzaykksyIl3bA7xMufo1F/MAvPPAg/MQX6GyP7wg6
YQof7iKaWxY9VriuyAiJUCoKKgaFfVTIaJCNn8Cd1j7zOgIlZ4awUWyFeATdswc5U9CXOTHga/V5
BoQZ6xKxygz7VTT4Fqe+2C5qzWXMSxYQOWXcGvDUZVt2Dm5LXcj5u20nG7MKctC4euBp+lF+Lzn4
dwZbPGHY1p8kwptWFASa1xBbQreeMITNE8K76MKcODUBBRPixu+40hlpJrgZD4rHaMK0mV65aLFk
vylj8Xr/72aW/wBa8mTrTb2/imgKcTa7BGAlUJfuvihUC7njVG+07Ff80Stn9d48tr5w+IEx+gcK
rc28yP2gRyjVa8Ond9vkDApNX7rTeIRFJ7pazcxBnpIVMckfwFpz9v/nxUTNJ++33Oem9xEnuifz
lJP4uDIFPABxcy6cfF9xiFMAkOu/dQ+C6CKpJqvBfSiYEPfYB3jBCJa6REES1Sl8AnExfJ8OjgvJ
gSvefVITfFftbpeEVnQ9zoBBc0ALadr0uscqOjNTfe0Ye3TWpqcnl35Ow1G4WcyALt7jWdw6RgrW
I5OMFWVx9dxPktwagxD9RkLQ+zaLJ2V1eDtEhUSSywrVlvXyxTmlzgeHmsOHT3e5OATiyEFHbJx9
n9u11zFulIhsXvzwO8amoU1NLPyMEtGpwuqqofL66pYF4kET9sbJgR3n/HnKKpLlOtHJ+SgnFn3L
HzJWw89NgA8h4pdUzVQg6wPb8xhcHZsXJmhg908HJ1L2XECC3wSUd+H/jkIGdNgS2KM5DdLsnh/N
yTKjZozjrjP6+G/OwrABbp3J6hYnYqzJ71QD/ckSjVpbg3FoJiY9qvTxJ3k7R8kf3Q2m8JBPZE+0
jGoCZYOd5xvdO0JabNpA6dKTb7SPN+YYg713beBDCkr/idiIU//Dlh3cMzM5M+sG10HBfDynLQXV
EfCPFYjWnL3ptVAsL6Kjvk1Q5aiBBGuIY1NpMqtBkzgC0z4thmp3Ov+wW1ByZ8KOCgJrTO4F4CDf
lVa2c0wZArMfIjbxLX4rp8QVuqbG5rMJd3aTV0pvAM7q+RGeQz1tDFBeEmU/JHMfnoYw0hNy3cNv
Zj+nVbzjhSp1Cs14Z2Fs0lWj3blg4lRmvUAweZesvewwipmIsG/K9uf1r/LH7iu6MWhAdhNiUTOs
tuXShJs/sB/iaYcmJE0vryy4EAt0f+fpM/DrDOxP+MNodHJQSAENEMKifpUfGM7m6w0l2bBh7hvS
H+BpCNEbfYavsO0HChhUw7I/su8NYzMx3IwMciwlp0s52ln4rDfPBVhrSeVI43Z+lmz4KMiEOguU
SfDdJbmVEY4V7h/ivhtwj7xFNNlbJVSHzXksrl46IFnLY2nNSuXRc5sPUK5b3Ack0wkuqpfuY03Z
F+uJH0hE0i5ebi9ws7XinvCp0ncqw1Vp2mM6UPk8l5EA00FzOaIiwMOPNpzI00xAg9tv6jD5NGtk
EavfXuRr8m10ktth1XPGTMqJ538R0pecP1a1HuEWb99MZmboAEiqrFau7gr/Kj0YInfF6yqJO3rY
u8RozdjxJhX7c4EpBhZDQ5/b1hjK508lfnH7MeWE0IEP6tZp5K/FauXDeZy224LtyuZXqXt72oCM
+Vq0e63LOYNjmCEotWwPDgXwydRpLW8FMKpSKVQjNqNXg1KQtKxh9PWZEvf0yLmOnYrNB82m7Ikn
LJFq1LipcYJk2YodWerC+e4L2vHp6t8io6GjLL5wQT/Nynoa5D72EniVx6cq0PMBtdLxjlL6sxbV
F4HdfkmlJA7xWPyGgxcUnb8f3IqQwF+CkJXSwakqtgx2b5KsiZuNRwaOGMt3EFDfufC7KUljZWic
UPp8x/UfIRht+9ErXYB8kZTL3VE2maFmGi391AiVIqb9l4FRptEh+fq61JcuoTEcDLJciEk9/lzc
v4bWFdwuzrWQHpinHNEJtXPTKUdt5W3cizdxCHStXOdYUiY4HJYUijfb6LbQ/4+AYK4WXGzYrx7T
Hs4dDML7Cx5gXfyMw0dO2oK/0l9zoJ8UUGwiOmyaUDXRcWchoNecNMRJfUprTmyR9A5MwSyKn1GY
eaw+cr+VqDBqkfsWyMWC6b+voA/TGvLNvfOf2qiGdpHAPZjQsctW4BPccNAjgyeLHZQoD0KE9U/T
Bp3ApmV1QH4vnQV/LKmYyMyvCtdDhgHlumK8w3b9sxv9/eQoBfGCnV/SK+fDPfSE7OFHq5Qut6kd
NRSq3zKNR/PAWT+AdAcCtigeWrwriDmotdKsgIE5V2le+RlWodQrHlz+UU7PM9yMo21HQc6Hevhe
PFUltpyBAfLqM5rDe/mgxXr7ODdTsNM3MoljXDd1LhyNvy2jl2vY/ipeUPLzf4lU/LEB/OrwizJg
hBHJpvWg/q1ZjMXIrdQfmJkpKP92diGWruXNlqIAkLjx2YsQcq4jB8vlMCNOjPZdpbZpZBXr7UCM
02LhgWTaPNisCN2AnFkHOz+17v7BkhKtAuZedxdc+9PKO3Gh8FuoxdkZpJoHlw7MjHijuZrEwyah
3FSRJEAo1DCohhbHAnkzufHDe3JxgxKUNo5CaAr2Upv0/cxYho1zVBwWfj/oMce6Law0T/BbmSvk
GiNGE/htqeTqMBaKSS58mKOzuvj0PWdnp+5X/+YQigC/gSTkZrtOTOR7AkaeQRAN2DN71aNFAycr
91eudS/USvP0fOyDKeiJwIFt6qkVwcgAaQWe8PwNC69F75L+rGtAK7uLv3+DiPyzTXSP1eyw8D+N
kWjSyUTkGQiB0HWOXMXap+qSOf1f8VmfwCPoi9Y4joNBNDdupQEfwNOzfGTo9bJnPG1wNRH262yX
j2ZTu2t4uIsmgvXOnTHk2/cASPemBiI6ek+40r+7JlB+vBr+NlTnPKykvdgYLfoQs41BfHlJ4CZe
+NWxK30YwRD6DnntJB3caJAM6Cb0xl7WogEBC/ujs73C26ERjEkLaXTmsADUQUxdfkstPf/ql71T
Q2/bO0kFxsq6LjnGpsG5XgrjKFNjw+1BMFIiEvGv4nyH0fA1lgEkct91IrWU7Ev8qfhZ9X2Ol5v4
mv0Fk6RUbxUfW9aGpf6fjZVzTKI/MxqCnhaN3ybvTpuYp8pQSl0FUAD6vo8xHtf2yGDhQNrbc/h+
JzimxLCi7+fMdCWdIqS/9Tf2PqMq6mA//wqcTZvtuKTgV9aUZUAZ9aO5IwaygYZI9qYVhqiG3R/V
yFdSnM5Q0DLO/LH8awCiF1uMZ2ri2F8g0S11Q6aDNLPonG0rqv2jU8hFGFbY9etme3c6f4RyiR3B
7+fhDd8bRQ/3euVSLA8X6UDb/1bbGM2SBFmhSVE0TwKI5EdVXm0CiOaNXx8zcyyJ4/ufMuG/hjU+
9y9HPbJdYJQffGbFxZiFhJgAIif3Id7rvrlpS1eeHZ0BesU3cYn5n+HsqIg4/+8jdjnXsBThUBdi
sJPR3ymDaFggmCpiqHvh+WtaxUi9xCNyBjeG5fYgXV81tPrZH8tAQGPxgHLghiCUlgXiwG25fUmB
pFpcgk9JOJjN9XXUqMEIIPkEzSFsL3Ef2bW3hfjKAW3XQCJGfxG0Ow8JByMCmXBwGk8fRIahi+p6
aSfQRU3IUu28jAHFFCYihJGApBhPvKAIQQfHgGwfRUTShK2RWeFM4p1DFaSJBCAVP5uRqZlKFlgc
KOOetIlI7dk14iYWxvuzeGx1OLJZym2nz4F/trPHKOWxW0TT5CKGhLb3utMP91Y72WtmrSur1iNa
78M7CM3M5rHXO3OG+g9scLIV/SMzw9Gn2DZs7xoZaV5IRX5aemJLEPb9KVjQKG0kk4TT3U8xqltc
sk52E5fsKaBMUxPg5W0AbG3+zmqbZaXjGzjptdKjCV7AhOeZ5UvImd1+Oxp+QSTB3dHXhQLfqoeM
xvUPgz8nm2USaSlRBw/suAKS8fLer+fy4Hn5rOXsPiq0DpyWMvzU4w9lx7CoRakOYFzGRjtUyFfq
C5NnX2iLKRzjzbyQw0I07v1ChsD1SB16B6TnuNH79AFdw/UWGJirmrb6V3Bw32s6/33cqU+TR1SL
WQXs9Xmdc/swcS/bndLeyMicZGeqKlU3dKvR2qqNZ9BAXalh8aMdL+q3Acnn7ZO5S4lcuMDv5fhQ
km+PoPmQQ+k0iTpJ2DUPwheMq+F/jGV6XEZr5w6rOnxRoNMTVgJS3ChMZ1Vs3H7i89yecyTEJrSw
8nT1S1Ba+Rhg7rLFNpQrrOJ8BauLEG78XKBnm8lMdtRuZ4SSGOJO/ujEvjMn6f9r9xKw9p1YeYyo
rP7ooAVVtUKK/ZB5/saffgXasg8UzwIVHJ9lFpYfmPThM9MV/6q734NwbbSZFaQfOC+STsfX099s
XI2RGG0ZSRr8sty/ULzXMMPIS78IU71gUJRq4vdWOTgjogUmQY5b83/UPUtNBv9+WlLrBamvoFaa
7ZXKzEgJghTfl++OVGRNQZMcZ6H5MdyuGhsLgdrbM5lSub9m3ZnuGpcYPa2EhifKmHrBFekVG90Q
TxrT7EqegaWywOZDMw/dt9IaHpptKAMyVfh8w90iFC8dOwcGBj1wi3Q0bqdoPgWRwBSONqN60rBv
NPDcBmSvoHAkkGCBPsF53BH0L2KxN4MC+XhcVTk0o32HHtQ4Jn018rtG3bb44o0n3G5EfYV70I6A
iFVNIVrphbiw3/UwyXf9GAuuI8BOeT+jqfgbYljuwI89sbJtX5oXoBZ9gZYF+GMb3eXsNAGoNzV1
TqNmwWjBN98XAdIjssCKIbUEEflpeXoxzRR62tatvHaXzyedzvLvhBUPdvmuUdg6nqLWKGCFe9sh
fybvqkAZVCYa1G0vzOWLIRK8z/31oP//zmlN8NgcAhSaUjJMVELjqWJMLFkCvIIRHlXQJt8fEQcz
bq6rk/sBeV9QrbBOI64lolDPjO6vChwYV6Npxp1ihmbQIk8VjU6LpimcmUG+w1aI/izVwW7KwsL4
PIhPbzblBo4htKq0J8dY9v9i3e/jtsaXHRf/gAbWKU1foHKqKlpdhQqlpmPpLI4TceMBS2rU+Hv1
IblU4xQ97GBBs9JC+nvFXxbvYeldefBfj5GUMECwLIzP7vSiM+f1swEGQ4/36aoKaF0tqiqGs7gt
Vt+9nXZ5FjWHSKDYgy72/akqW9gqds7E83NR4n/BCgIdxuC8ygK4eAU1MYInCXHwr/cTcu8x30EM
NCxHJUKRbw/AtDlww+WPR18q+uYwkOhqIZ4vHQyshne1cSfqLIpdQ071t6z5dbAPpLHTo1zZA8Qw
s1FwEsQL2jSp3sRom3xeaoZBrF1cRWO2u5OVZ8MU2XYgDVN5Drd7SaUf+S8PVoEjcQd8r4iTwSUe
+ufkYZbdGXEgYF0gco8a8Y+7Ii3OB9UJzEyveZ1RqwxLouEzCLSKyOJcEtg95V+q1Fhd4q2Z9yXj
Qod81udjD9OkxDvVk4nHq+8J64Z9l3KzmkaKmoZP0uuEDU6TXfNyKO4mzf5bklkTmKAZ3/gut9ix
4ivt4YN667XPlvZryhrkaggZ1CKFvhiubHpy+ErBqJHql+RyUx1De+5GM9W2wprg8YHlzPUO584+
4DfXdBhb8VNtjxHTUpJpkkJThaD4zFb0xj28vgBDL6KVuna4UiXZwzuYR5ND9pEbyFPxrf5bSIlF
LUroV1heFDf3MpN3rVN5PYQ1cuKkA4p4gr8MktS3m2hY7XWtT1jja9jYtB/cLOak9+oJoDYUnUdd
+z1IKyrA3SIJVG7rLt9eaab7w8zLRPh1izDK+XsD/qRFhLollcAQ3XTbDBUL6MullNjlmeglUJDZ
N37sSdrhIJQptCUStC4Syl2gGfo4iE1bCAwPOQXGaUutPQKVOxbX2KISrMbQ9KjwsqOig0t4J4NX
p6/KN45djXoFFRc0bPHJLM4c62YIJvjKCktfgdC/aMDv9DZBsKr69DtAY2AWEjo//VRrmB1n77HE
v12D4ma9tgGqDjnicEo4teHjmWGXQ3HamMFMOYsmPx3oR7Xo0pukl7oxIPmftpHin5GmjF6lLj4n
siUxzyPbJRenbHXelXEqYkX9iv7g5h8SkhwtIxJpFqpibIxtUpH2ymiEoWHVsobtaTkEyDwq/lxn
5mMk2ULIkt+eBPbEhGoOh0eVNsAwzkBXHj64ZMILjSsPWMByH7JueFWssJR6QzdRm/Xv0znrEUWe
tXVpgh7AN2WLRoHpPr/Iz2Cm2+3/MHjglAG3qAyXpXXpF4+1tMq7X+Dh7jsh6MRskcZl+gQ34vup
40tfrTjxUPZX1K8knkRmq4o36Sqet7JxPQGCA/eVx2uEjoDAEI7vo0P8pGN2Cf34kdjC6xiwlMhM
tv68Dym0NMmfQu6VYru5S8VY7A7Wmzb9d1xc/Y1OfKbJRB/F0izYG8p23c33vx+ot1YIAVkQJCU4
Yr6qunS4I/xERzgzaSD8YFbd2ZzzND/vCcf8aGOgvZenixJlSlIsdRjoNA/Ykg9FbjoHxn5ggb7d
vDMJfKv0UsAHpS4zMT3OMflaWI6LYaJzlAi5M4J47+RtNCIaVg8mWDHgOOJ7wjNuDfcvpDHQHSLv
LofA2wNdHMDMMkDzF4LXUjiPfxLvdKUDW8GfmdnfyLlxE9r+A8Ynjwv9WVkDm+Zhea+H1b4XU6wO
ebFpoWJIAP9X/rJV5r1uf1FFzIheO0VgT63Q/tqEc0epPva0eCnAxR7RBF8xCA+ytFVKAMxWhkVC
knAFfYNSM/KvMkYpqaC6vTYeHfCH5t5aSnELKOfp8BJPNhjxqxcU9vyso2qoKyrfvD8QeYjs+6ky
Ou9iahbr1lc2/Z1aG27R9wl9j4oF7eb6pGrY4bebXMGjuLxlWcaSrEOghuE+HfHINXSLDTWxIOcv
R2GFvS546TOiz1zQ6s3icHggwQ0cvrbHDRjpcxQ8rLtqU85ZyOV6cXQ0ISYF4UyPMw3INiKf38eU
NwKBFbzlvNYoVfgo+dVb1It+oHOra3o8wh+b2Pu92gvETwS97N7ALJpeQU0i3puxkVXNH1pezs4A
/0eoK4gqUZK87dzsykyBvR5MeW3vBtUb+xB4DkmXnzuvX+HE2u5Y00VfzPppv3wBe6P3wuSxSo+V
KVehsvQljK9tVhMdRfC/r+oMmLGY7qAanKX9Y2Sy3tkho7sdlC0mpGgdECGijzyKv+kGXEsWEOIQ
slA7cJyxWGRkEQyLzTn22gcr4PuEx0prZ/Q29q0Qd2P24wxJozlsYzaNI7eeRQe19FU/oMu+xFpY
VtpnxeZqVpGikZy6ooB9cbBnGJx//4dYSmtCvKa7ElUZ7d6nHnCdHT15s6QZqy89YB6GJTjOb46n
QsR9l6kkTig4Qf8Zw6djT99i+OLEZ185BuDZOjGktgwteNXj08beJiZqdtoyd6hKv/YvF/ogpdLn
Cn2NRzRjoUbYqXtgD0bmUk/KE5UxnupWcOSSMpbui+5ENDYU1twqhcD1HE1+vaisn0l8gNRNfaK7
HPHD6R0rRzKQ5k9rp558uxMsSKcshvz2T+7etm58c8sZNutwzkZdYLUSj491A4NvZUbSXzoJZYPF
k8PqV214gxHhu1paoP6UCNmJP4hHVodAHn9BKbsfZh6NyLJRjABW3f9biTS1Pd0bl5d1I620o1w2
XQngOC5qKtrUqvYQOthATC7q2IP+Xq6YHL0DxOQN536tE2RB+iB7jixmr9fj29XY++Ld0+5UgFRu
m4PZ7fWjGFCUyREHkq9whhedmFX4Cc0hsuobjbgysZCbqoZPJOqd8S/oqxGLNt/wUGT8dWbhn5gi
fqfXFU4zQuWUqQXXAs/hvhP81qI6683AAiNZ5O7PsJVDZWZKrYn5oz5JuW2PteO4IGmTzmlUKSH1
667p/6p4Daccq3LWSy5dHpRnnC2Jv88l2YxnReWS6GQN0YsDtjRNLEIb+MZOwKTBBKNiuESmn/9F
L6sZBi1Q8eyrrx+2Gln8wcIP4W5ALAN75QwZyF4iOIu1fsyeh0FBOpL/aXTzEoHb3M82/On67oho
6+UpsywgKSg+Z8m48b+Cc/VrTvhlstRGjbehixPC5ZZo4i8D41Dt1+uzgOKMHgkyqYFbE7LisNtF
Cpv0Nbor13Tu6fP3Dh+1YenuBhLQVQAmoRUqj1NBB/nR8rJCb1JsXtCp4+az2Fl1BDtOObjrBraU
b3hp7yAXjgnwbq76rVjWHvuyevCTgDu02w5P6fobkYX+PjHROTj6EmcCg1RojrArF/lva9ikuL/d
efM83ph7EPGCwjHo5zQEifursi+23MR/9rNvchCsXIiplzgfQI6W0WfyVKb0xwOX1xV9Nvf7gjq2
7a5/h08CRC26JtHBT7Y5BxlgDXO5Ey9aWeuvKPeAl9F3Vy6wTMdaZZn99BOH3pJk6MXzmWWdSYwf
ZmwV6ta86NlOXyTDvGo26BZFVLxm0Ax9nyIXDqh5/LobHuJZU0Osep4KMpaAOwgjmhoEpTmI0K7b
+65WfCSESvfpbXCXkwSdUMd7uNHOhN+p8HRyiJnry3XuAmkHq3g8gr4hS9Zqe5vEfQRRrQS0O5Hy
Dq8g+ODTq7t5r2ZMm3CFkjaEwUa5zLdHbkEBOt948lPimtK2fZrUFRSnMaVIzqHFxOgjgoVGol6/
NbUHTlrJq0dGcACbWTEfRpP/4j/IMG1CLdWpyP6QBY4qZIvWjfPboj/lveNM/d23m5Iqu86F3ajY
DzRBWbEIDvR+KfJSE8SgGgC5SqhKzc/gnFyvD7GeYMh34nQB7OBPU9Os6XNi7nsQRla1kU6dRkeG
alAcMt8lK2+MKxu8r8WBf3IW/2+rcI66NRHOpgkP/ifwPy8hOc7jlRKyqllp8x8LzwT/PgkWQh3E
TUf9yQMblYr3xxpo2hJpqW5+QyMiAElo8JC90AxdWeiB+j3nS6P6n5pOy9Crir63LfL7Y+swIN5p
3fnTFaBEqO1zQMiw4LCBJabxrIksVaHV+miATWadbEUZAg/V4n6SJL1S/B4yEOUjAuYHqZnCeIl5
ttBJheGqR88KCl+AeuXW/3gL4MdtQCaJZqd5oX0tifNsucbygNCf6ptM0j/aH2MQKt0NcpQk9oGo
Hvkzc2TeCWyVu4phhWKp4ndhSLEY8RCHgWr+r+EOd6LwFW2k0SUeOVmpRbOAq55ZKdBQDECpYizf
l4QErrb2mUugVgDUDUl4o/eN7kIDeLqlzhMHmoSEHH5TIQTIbWoL3HDGAV1fDfXXXsUmt9uJO/Nn
+P57dPGbFTR7L6y5FDqvTkaI73qMP0Up3AeGGikMa53nqEg/yxvGVsM0ApQqQyinq+Lcmt7AdY/F
NXXgbW+//go2qNBBrDie/59cA+a24Gs1xkBLISaUfEyzPYGBfG5PR8w/Ga7Cki1NiizTze1UzOpl
capDhudnQygf+IWHZYzlZwRNxmGJwG6gND9ipHLRXmGOIP6PLXm+Utlwjav6x1eC/C2guav3OdAz
LXrsI8lQxGm+KZR1a2enxxC4oBEGUAMY8OpEf5NOUxE5udn2CnpPgw1WPKVaX+1IzUDMBN8MEbHM
I8ziz2/94kPIbtGvSNdtgJE2j0NLzYofPuAEIJM6nTPnyD4ZlpGd0Z1k1xh7GJpNyvdd57shExyk
tkB0OmzDzdoRTAmwUtQEoBIFDD6CKcIZRXQG6Zt/P+cz0UFU0eZsNxgPZRNL2AyUfN9Hj3Eo17au
RPclZlxN4VnOOSKsQZlN0FrtBkY+RoHDRK7Oc8ENw+p79y+u9vb7aexeFWvzjaSTQBOZJwf/4Eus
XMJPERc60+lV2MbdgZVv+lXUBqmFQzB1UHYnbhhaUiYbTzhysiTgD0KGrD0MfV/OkNWwEth1db1k
FNjCueCab4oqPeG/aJvoDMXG7eisEd5FSzQaNg2Oqe9ZjOfWk+e1dxFgKkAjSFABsKMdKErb16Ws
+HAxP8m+wB3+ZkcYPIHIwB/blN/1rnnjLdQCuTp/13bDnO4POtM2bqBm5ZtnWjoGM2PGxNXAg4Iz
lsHquxPyFPs3arwF5Qrc243/4MLnU7QWBeY7Lc5RKdIKiSc9bVVxWmO8jmFnXsxYB5lRWUjQxqjp
D2DlH5at25U9m8IQt02DVj/wIpgn69Mtx8xzTlzoRaxaGwLTJoa8HG4Vy/keSWnk7RpNnqoyZ7cm
1FIMIgd01Y6IOdXPaPIFlE50PPUohJ31a9ZXIGSb7tSTLq24vkXi6ZwDjSnM0FRb4ILJp4OSeumA
wu5nzjyhhJUBJhfmu2nYvPwypwEcxxcoz6Y6s/MQn7dvfpm0LMYaCQ/e3wRqY9eDCcIJYQLalwnj
/5aMXZr5Qx0DaHlakScK5UuQ11fZ4dqGUP6U15fi8peqpRtwXUG+HqzNeB0bI9pWKLdY2+SRpezt
TTu1uBRkcxqFWrjvfIq5AEDnONGrCIRStg+DF3UgWN47fx0Itw5e4VUnNnRvbPJv8NEKKvrXfNSt
gtkHo0KoFEQ9H5TtKDOSVMqhXKGyks+hucTUSFimZbQhb+usmlkdjTxkxRwyr/U4DVKS5TJITVNz
neg2vl/0aJuvqNAO8T3qQeuic7ipkGf4n+dxtIqnrOVXvBDJhhqR3L+1oFsLtoNjoELGZ4kk5rG3
+FwProAvkAeitn6KY3mjCtQI4gJdf9ZUOu9pkXuaiIzSmyZUk/5X+3HE5mxVwdVw89fFQFeRtTjN
153L8xU28LDGG27Mrp38VPmdE+6YykKStP/EbiANeTIziIugwb17tghqt/kA/1cueivSFre8/tZ9
9wvhypssTSCFVCBn6WHJZ/IaxmvYZHji9gECFZjW35kJYxS5j/pSJ+kbQF0DmqorJqByaye5BbIi
1oTyL9n5uUeAlYbFAzDhBsxxJ9vxkU62rQcYZNtxpdFlwH/Wa1n+MhCwPqqzFY3WWmB1vF6zdjg5
rAytNR4yWJWIJDkTRJX2ILpMRryBPZe5CZ9psjKwX6ZwBPDX1RAEQAqKWh07dbzfdJh6qJmENHwV
Mr8MrMO8pMG27BIskMCttq8MajMQcDsYW3wOacuojFqljy81n9i99HpYBWK0jECr77rDS90IYEIP
X0L6eTdbHSqM90E2jvzsspvjRXmYrkFVhHmaYM6s7T8kiD1F5OtLnAZgLplwgUADe02uglWGsSgm
bVjzWzXWRgVyjHaVdmI8n0+KRS+eFzca5QPUZTrX8KOeSgDzyG0r4Qlja5aTWqKmaesTHJxYgLaJ
+vGChepTUTaAAQg1abkyxWMzJgs4oPJjz8aesH1/WndKGe/PA13YKoV3YRQ7Rg08AET7eaH6hNBk
KLM/0ePfz/n97FoL5gASj0MuHcDTL0T962F3ri1S5bDUDt07oLnHnrwqbVBivUaysHL8E0CUhGBy
Qyja0rwhJ04TYhfCnTp59BgRtXbZyBcb9aiA1FAgSlf2Fh5IuIRXCIAp/SjMs82XUE/FOj9HBYyw
+RMmyNaF598eaZT2mTWHEc/Bjx9riLz34+adHPzSn/znRHC59q+0rptjh1jmI9aGp4yR9t44693E
poDqyinG32MgekehbhEC0LXqnQP3VJiqXUtluydFScOrI/wK3GYISF9l9Qufgo3YxxMdSd5I3uco
s3TWOnrGfTlwyfHg1xlcMsHVl3BgjikI+Owh2hQ9E9IKISlPCAaPEfeO4jjiQBDCMS9+WPReYMrP
SZ7e6Ls3TnDQ0SP0d4yXTr3pWjzT0l18i+hBeu23hrCTYZlFTQ6mDsVas3OHLFrUKPityj6skEkh
kAt9HP9pr2v71nWEqBaD/M0TfsY61dy+r1c0/J2qKMoxdqHKvl4nkSITgtsfUw7pKLhChIVFlzQu
/fPS0jYl8nFw0O29Bqcx2kx5YnxJszbMv33XEsarWN9/KlHfZp4aGFijmyDD7F2VElKbP6A26GNO
XBwtvhkcVUJebQp60UYrJWTrQEjo1oNoqx9bOGSr6+luAjTCPDKDQVB/AwnGNdfVTyQjt3/UhTfo
r7nbMI4rs0IrfkfqBhxKUUNMLBYhO+wn8/kboKMqMWu2cz/ZgsdTf6mJSeEvTOZ4hBQ1+C5jZwm/
a15jZghvEhB4Z/tVuhOX3qO2Osa13qZnneADTWOXhHUaPIWjNBS5Lp9PocGJmEvzFI5587wPGSvt
hFQMe7PoQVK6T7UwN8738IXUEbACnbFR7EWTjJC0cjdy9p65KksKf34UTg8NMw994MseY0zSDNi5
UqwicJppjhchGi/uZz8SztxbtTYUei8G1PYuPHr/TenyK0wVYKx1fnjp9t0BeXFPdR5puCAF5Xrz
jrt5bVSV6ecCjn7UfYgr/17eFRcjodYmp7SX36AmN+XG8sH7rr2FjPYY4GXNOu9HwYE2/AMNRfBf
G3K5ny2i5+sqMB9KFZ76ri1L6eeGr4urNQcj9igCXW9uNqOH/im+WPDscEf17DugNwjNGPlCCNFN
7Bh2qyrz/KoKOG0e3BNGhvr6wn53wfyEoqsG4A9E3wikfygfrgBeExWHznkyKonG34Cwwp39oPmO
b8l7FreHaUmO+giIjudxwB/us7U14S1n08px50+VLGU+bBNFmNO8X4GrAfb7dHC+1UoPSFkkV5EJ
tucvtUgVrLt20M6wQJP3bPHS8u8KzpAwNl8rpt7FooaT/M+mrSEG95qPAnI7Wqdf5YB/DhQVZCGm
rWTLehDhlj7T7yWFZcWeZnP90QrK5Vcx/wSlYKsIzh3IMrvf+NFK4IdiGEjI7WbPBpZcICoqJH9T
ubLrdmxX5IOFFu8BMBKqUpSGlsQUHgwb+BwDuf4wLmaoFWRUtmk72+Evms2bkmbLAz7xz0q6wUay
4G3jYF6SuDSTn/cM0j6yLYNvweWgQKnQgfYc2AkW5Sv57q21pai8znpCem8WLcYbBdkmLxa52dd1
zbZrlfY9hVYOB3wbQzd9lBDD5E+K4POx7BhyVlBBp/TmLB33gON3eACWu52FzG4vQBCMirb50bdT
p8VlX4VXqwR47h9qCZOeai0sBshnWb/Uh3AkLiyHcg5rc4Iws2CpRzfYdevL9VHRe9E1PRab32a9
46L8izGjMnRP9F5WX6JSbO459/p8ZcjS32hQ7UH30GksiPP5+KI6nF1PXtL3KQN6DeIKvtgk0et9
2eXchg6MEdcfALBOhvZZozcLSC+bvU2UIC0UrQlLxgEXUl7H+eAItnTl8uotgLdiwEN86xJKI9DF
mTG5pSfm9pKkf36mL1XdF4Z68oZcJkhL/xPxlvphI49oR1fbjL12DxC+I/OOH6Cu8CG/XptKFysq
i/CEWYfmJTl4ac8eNpt6sKUkEei3RdTtvEB19qgV2Eq+VUbHrP6OWYHRpisVP/JV19iyYEHQcka8
vtvcES1PXoZ2kK3JNYajpfsP6tpT318oNS0llw0FYQ6J5+D0EO9WTZ4xnRACrmqSzFvduuPZHrGw
idIVpq+6AWk+Di/fm00vEiZ2xvVlQPzXIkePpf6F9kwD+3fuEG6f4NmJmDdZfukbk8PXRZBmzhjJ
XIqq/+uTJKH8mN1uEpCCsH2itpiMNPRAxTEjleUqddJIbwo8NfRdsDCAQDn8MMhfueznA7FKIj7+
NV6vv2iHkS7J7WcRItXBNFPgE/+/IDkjB/B4NN6duG6o8RzGDJiQOi8vrme3Fw8fMGIx0Jm2oHTA
LvnubC63CSI6H2c2QC+QRv+r84JEkXNmdKC2rtZb9RXhnWJ7VhskUPlSH1k5GKztLzgiaVP1Ilcp
Aa6watCwYjPLWIuGw/ey//ZL36v1cIm9iu1hy5TyPgf7tGS5lbCVHdEVSDLGoawIH5gKpmHUy5bv
JaTzpNWbfDvU5BeDJNML6NtJA934jkb9QYnJ+liHfDNCpls8iecYM4WgeejJJi22M63grQBDrBK2
r308zBBTS6B6coLDTs84V+pT8AeUwZlPh4C7LFY0+w5k7tQtVrixo7Ow9ziHeKLKqlbbcWp45oGd
ZPBlqePfu5j1QoA0nxfobopgFVwRPfnzMlzAQ8WKixay5YlMXhYEZsowvTuEbGYByFtDEzqZ+HCr
8lCJRM9qFdkmpA3/knHt0vWD2xUXrUer3RPa2PkmWgs7oZSRuiWEDJ0Ig8U82oDr010VKwnggrzq
+HK0eVdCCK8ZeyUoR73EQeioooo9aBwO0dGmDIGLJB3lznqNaZvm+w6mpNaCqaapxNnf12q5opkQ
i7omTbyRDrMKHKxK5Bh3JDuziT9oBMxrT13plN752IbPmHTkvIbrm8kk8SafWxmd03gOO6c55YyV
YVx+QWQ+cE/xrOYEiCI+A6K4MBislwMDr+hemXf8EQnoXJ66j0eSj32uuMk6BCkqgHsaSpbA+Qsr
IF6KhOR7PbqP36svQn5iJkDUzCzgi2dEfWSn8vLhUCENyBFDJxMfwikK6WGVJdgT9L5y5c5GRMfY
4d9tqsFp+X64iqAexTJTHUkDKrCIfMllvpYPd5hgj+k27Aj9/JwPC6+PPoq/0Kv9aXCHCiSIuEXW
SD0UTI1wI/1qx597k02AuN4a69KcTZuXiLG5K1/obldTykAzZz6ApMgSbXvtbCZDhwTPQy/f+J2V
zL4h6LhVnDV5RqkSExdR8G7KqK9j6Dof3fEKj8yBaBre0VDFlZNFlO46UMJjn+HmuKaj9QSaL0F+
WRlzgYpSCrOWxxo60RIaR7XIGdwa1EsnU1Ip/IgTQWh+IMO2KsjYL2V/wN12uQL2anFeDCIjjbdf
gw9Bdwn5GVhLjB/embitIKIWuenOmnsiGFkhMts0plozqCR25oaAUxEDxODkyEbw8Owe0Nk1Mom2
ARSW9Tl9s58K9G425bP+d3GVVkAEsivnPyqsemb0VanDm4t3w2Vj7IY07Vq3uEUs091N506gPvek
OLE8yx2oV0ybxZpL3FbXMooj5rJ6hKllAdnF06K0hEL1EANfNrq3vN7NeloOOnKx2hHnhvNMZ3kg
hk9c8S3S3G0cBci1bRDx1zNYnVxEz1ITIzkCu3DM5o3iGUM8aOLMH64m+m32fhkEzWT11mZMJVus
u6XAfXEN07/Eo1yAUGLvKpnSQFscDf2cCucQAvlO7WGjCLP4MQvJO/txeqgjEEC9hSNd+dGJzESu
9fjZOqkip4F5/CYtTkMqLpf+23g1HxlbvKDDQ+0gWxxt3LPAYTp6EHWbYTt6PPCDJwbYQLieKPiB
MRzMSzRNTKq8GJuL7IfnPcPKiqeREcoAoGT3qrvQ31ICjPFKK9Po7RmUmlZy9h1rOUvL3qCcmZd1
k3vQ16+ctfNdEfdxGjW2cVfHNstdwfrapnGmmTtnBpYO8/Y56MPg87fXZ2iMKYG5ZRt0eVqwetQR
NSkyXq1h+ReYoPuIg6W1BqUChxQ1CpaznZ60wT5picszmoVTohHNGK4PxE+02WKynMkl74yDzT4/
pD5B3+LkvRX/3skHI/j1G1YMJ40jbzhC/SBIgtC3SfiV3CN5RYC0UMlnWQL3mgDl0nSCSpussWBB
kEIZn6yd4bpsfOg3Sj9v80QLLQWuCiv63IGT1mgWCA6d8pP/7TdU3d8moHO9uE3WFV7dOF2ipnLi
SRqVky2p92hzpbNqqcoGLe8ds7ErNtCSbdPD1O2C+cUruwVtbVR8W/1Nzd8jcwhI5spzRSIeVten
6sC6XkFnpCvOKaO8j0XpUrFyLD89eNPeFcYDX9MqNH9HbJjW8lRZfk7JpgXElsiIzMXKRBKMw9bP
rudejJNEXB45oEEEHpfLkQdVXnRM4qU/WTSj+2uJS2okvAkqTm1qirAMe6dF49+yQMzQGVYnNSH3
/yNxRHzWxZnJ+nX88adAvoXZVlKE/BMyxpO4kNI7KT+pQxfJCol4VebIXHome3g98hybV4DqT8uC
9WlP5Jfx8DBaY63WdinFZN+eDSnFYEaMqLh0bmtd7l7kAvvLY3+Y5VnWwkrMMeCkektIn7u7OYMT
y0+LyfES5eYyDzWGQeaosg3YAzwnXHgpXO56HIjn1sS1pnM8fc4RqjsrVupKqYcRnax6H6C6Ag8b
ai/3dZFkTl628t2ZIoR/whr6BWzoP0TecWa4HRxcjQddOUxIY93oRv40v2Zce2W8deVw+imcliDq
4vXvJOh66d6iJWdAcw+XY7ALVeEdMLZ8+mjQHGozCydUcKIthbBsCEmTbNmUos7YsdiK8z2wYDMZ
gBWIFMrbOL7sNa+guaFHxtP4whhY6du572Q5gLsnlFbcZ98YiMPuQlLK82sbpwTUZIGkuW5KhuR2
gl71EGN+9yA+z4leGyNNUqkYvuaRfN36iQ8DBEWAmMtm9vihsc7JcSm6TDhM2J1LCqewxTPPBolH
hgMREhcHimAM3APLqdQKAw4+OTX7Jq1KjJ5khvppX7UT1JHNAUw5UedAyOjj6krsQSkNgBsw3xh7
QIjLn7oih9AEPBll107x3V2Ertut6wPa1fdv86QaKNFR4H1hjC6YP3hK5AvkzUzWxH6WE98P7VJT
nhEU4xTqmctHh/fNOYBaauDWdVM+nGNq6xCH26Tn70Tj135uwxFp9C8sCqBRFYJYu1/VyulQZWAe
6pkUr3w3wf//3WOXBUtC+M6+8Rkmr3YpJL+aDzys/xe0B2oT0ev1xtnNhG2Z3Cj9QqyrPmAJIzKg
5GMCgAcgd3ruZ3XMzR6Ay8Psf/K56iAPXIUciHYvFyU/vSnLGH+gJ0iGaHloYTxLjonpSsdct3dZ
RqKpblmN593uKAQKwELPTvkKpY2tUdCPTR6YQxn4Od2YzPQa50DrTBr5SWRqHyv9i9G9owPw09QV
UYNKNugLH+pDE2NN+Df9I5WjG9K+qxN6e7V87q5728T57i3VCD5aMixytofpktN/71MwriEDP7zQ
D3g+SYEeDeXnHVyPzRus2wfjEOsfzl1e4bzrowMZ4ud4dYxMo7/80hgqqTmGhLaANkNmS6UOjdKS
Ovayodzlrsgs30YjSGMeNR5ERZdg/G64orgWjJOjCjOjzYqxGu3RGr9wX58Yy007TvgPsH9R3HHb
48AXHceUtFhrGhrCoSyKcSHoca8UDf7uzfkaaY/VMxWFl6ZMSgKZ5Lse7BCx4Bekwig3+d048F34
2sh1ywThQliylPP3PUfSeXDLrl8bCo2a7pcitK8nu0mF7OrkMqMSN15z8rNX0ZOqD4GvnDGt06cd
k7y+B6O6WSkukmwytNbh4sH1lGGCQVirmnj0c0n7HmdGQZNQ5Jo5PYIMBWNzwJsg6cb+dzLTNA7e
gLlYpkj2RBKi0GDk+15vSOIJfITpzw2qFqkDtO/Y+okTDz4aaA5O6AYUnofF+tgso0TNNNJlWNnx
cZm3gu3lHkid8UQbjO2rLInqIqexzgFBtc8+lwjiZAkRpbE3dmIUHxQInUmqi5C6LUCPHf8nzURB
vLMYQH1PpqzY846lBKYG9t0W8zxfKbX3fLirp0yUAK/Dq7Fipv8fk/ansQh2TMfqlNgKuwyp+87M
IAhktCQxa6f1J7RbmFWThMIcJc66onXEAI5HX1h+MMU7Py/w78eRD9w0EXfjGiMlThdlMm169mFx
zTHn/c/i+AgrOiMB3UjGFRwBkZ9tyaFJTxHPGxFDuie2DJ6iP8IVdUtAsEkQqUaIbSVLpaa0Q1RE
wWjeh4TgOkgFtvF5qWjKQtiVLoh+k2PKANCQCqG3itzi97wJaKQfA3R24EzU+EuxsjK1iozd/3WH
p3glZ3CIuKVcgubwjH1BDCSQd+sEeFSY0Ya/JWNwi+A13BAge3srrZ9SAgqEOrgnu2YsnxU0zXrb
AlVP0UpC4NQy9YxaNoTAaVUVhzZAvsk6o12jcd+jyEUfe3YTVvM6+2GUeNh6ERIRU1BNbjpop4eK
QZXI6FE4SP/SBqgJ3pqiiKIw2auZPV5cnToolIl2y/+xh59lyFMSD9hcnuVUAuWqeexZ4IMGj1qq
R1gaclH1R5oXVwyGd+fFrZX8PT85DcUw7OdoVRicjDRdvm3Bj2WqiiDbIq6OBMs1wE9/xxKcSX4h
q8411se655uHON511BVsfaHWRtB2ATZdXIMRQeobBcjYxArBhNih1jBqRqvH+4FbqbH3UMdBdT0/
gaoN3NTjkA4v/muNg1v1C+gH5GUENYdWm3c0SyNlW3bQtumHFhXff0/9Lc3+SWcoosTn/eF/v5ZA
egTNKxiFGTX23i9ezXPbSKKBSM/A4AOjATnDlQ6qkrteXv8O937ao4lQKT4wRK/0fsL9et3pdmGt
QgTkI7U4d52y1GPYtXYL2q0XdcrIZe7uXPprWgMx29hA27VE/rixUSWiFRd/+Ce4QeJIvq7Ho4Tk
GbDCfdkSM8MeVJHC6hxMLUtDn7Tw4s4AZ6CY8FOupG4A/g8JzyzG6SXvwM2u9gPeYmsmEQGi/HVp
qYmdjdMTzvdNV4P5PK9HxqO+Wx1iSH7DbncBm8J6WmFQfZ/sDIBJbCbk9owdtW3uLqt+A7/rX0gt
OoPeSIU+CF8XUbanI04JqSVz7HDjLPwUJxUF7lKz4khM7JPBKfleSefOU38Zw3ydW1jPZhdmv9wt
zbq1dAnZgamjCQIkMm4orJLRM4hXY62irxJkdyguL+2YrGIlwUJJ/SFejMlELDfJuOTuH6CopmUF
r4touuTTbFwk+NVvXRKV0r0fDMVGpjmL1XAM6gj8iB3bb6/zZUEmoYDwqsqh+P6rctIU/0cJrj54
TKAMPjGZAJhmQ7NuOMhG2+Pnv1EgtieyNSlHRGymvjT5oDWG2ODMYFPHRCVw0BPS3kYXASY8RRXt
YzzFUpPOeUBxqN0Um/kHpdhrNkIvubNfBDcONtDVI2hd/I9PUjf0Q3W1CiPiSfk1JCjm24Vxfe1z
+BaxG/3mYUFcArthTx53Ahar+6XGpmq0dpWkKGkD5WoQNQUYsuPRoG0NiHHm93Yzqo9Ua2DX5OuY
wJdLwSV2dozJAc6C+xk9hRZHqesZPw80arpMZTtFcjR9drzfKdhmdgKOnWck7AvcNuQRw8yaHg1U
5GdmabUhUBxKQUcylcNpd5CKUvuFPKeAvaZzcSI3lhlhVd8k1mxd0JjSH7j34yA+BKCe1LK9jfBl
7aUlYj5swtXfF9EWHqW/GG8aOzbyok2kpfCff1txQQnEYwVct1ya9UvDF9UnEch5kW+O6zTjH3jv
dR4cbJtlSlQP0C1xc1MzoEN5umZVoRocdno8pKLQP3BncvoR+W1GSj/5E4wtE1bI7QOI6pMaGrvs
M2iJJsuv60Ci4ntP2+ThxmdKXgwbhMSSRa8mVHMj5pT3jL7mMXt7A2uFo9NGSppIDMaXGo95OzyU
KFEhxuQ2towSEonorxAJLcCzXq1+YG53cs0k9xR3aeHaXRA+qSCM0z+Lx6UgCV6+tUjHZxgaazZ9
0+MSqY3i/ziBTpMfvK9MIvGDnlmXJC1ME7Uad/KpGge5BfnkP5+y1YgVIq1tQoTZYFO0gVfAMYGv
vN5tWlSXrCDEYybdGTVPqZI+hhORgo0jzCd05IhibOz2ZMnMMeeY1eTZQ0oehEN5q5daYUdw5O0S
HvQ6+hhZPyLuBjJVRUtLhb1nAvKWnoO7MmZzqE22S6/u9Je7PJtn4LMBJHZP4BPJ00xjr/ww6hQY
Ekkom2LEURvWrG+dhrDtMoKJU6yXlBQxtVxf/PA6fwwqRqG0R6tpW7wAUzYVwxUYtMv7wh0jgLJ/
iYjuliBZaSyblxz1B7kOPWygdPFZHaEl4v1VZ8XGwCGNPMY1V50KM3AnECFuCIqlo3WlRkLXvvdc
eug2UQxLti8+rHEfOEsVh4xrcDteidIWERC9Qi3R8UAe3yU7Bo1v7SSQmuEK8Ooaw2vYYL92nY9P
fSxzqMpfxP7yuTD9A8pa2Sx79NZCfE6VYmvnwSqPgWpbKi+aJz1HXxTiY5N5OJi1JqNsGu/fxeTo
65tLAWSvl7+ekRFEg5GeYaSEzMwnomG13FD/9JS43+wi1DYy08ulDMSPegB+fNyBJVC6JI8o+vp/
J/y+Dc5sZBdQjCNPaOmFVOOWW1t/q9Di3aLZ6+QhaZnbYNDNrgUMdgv61k6IMES+cRhWS6ac+IHB
wo7EHce9krIH7QaYg4prttHL9q5v+7cvzkXacA1z2Z3ZMwQDL4t6lITc9RKUtoQ3ynKrYjiM21Gi
pKMViq1l5w92M7lelG79mRmw3YpVGikBa6z+WFbodmKQhk86NOfJBmUnm8izct8i8Za0hko7pulh
/OE4rIsm9mk38/VDGK2EN/G4SzmzyQy+wtiAHTG+9UToyqzQy/ys6fofe+WcuyulbrrK0bRfhWrq
hYB4kwSScvF6G1hfIN08Q2sinp6uyrx0Ssjt0nrDF5J4rOccVAAtY9ONu9A7uTMwuFxHTZgPWtzP
xa0PEonKS7ZvmY90lobt9vt28tgDq/I8dpwi+XL7mfRis4M/pkO7tQssELwkDED0dKklkKOw5VxR
/xyp6umKlOfvI2r4TVzbVYUrUwJnOmuM6xNS4qDLWrdrpFoikFqiiyuwexI5YukEUk3qVFSlb6ot
VhuXfdOWoX17UtHigZ2LPKk+ShKZQg8u2I/w5EYD63cvdCQWPeZXKLjtX65PtAud60bx7SBM7mZy
47AR5ovFvl5pfbtd5G66ZeNW9m5MO6bsLxbvH4EXqMvTZfou6HcHMbf54JNOWCpFOlRC3EZgoN+v
T9QEml4C6ZZP37dAOvuArfiTrDX3cm0no6cbbYHsGfPsxhmEX7IH0vZ/NUQYNnbwiA/JEtpsuYiT
gpluvuq1TJgFZHTJFgCiQqMZb9jxURpYeXrqmoUyOPfpqMXRCp1HUSwwdhxMMdyzpvngKcyXlKQs
aOlomp2NhAZl+8wIxbx0WtuaFqFHEeINX35DM5LjkG4L4e05eiDHIsrNV2TUziNN8aqBnmPmn5h0
NGVwBdLqrw6J8LbzOUebDeqsue4Qc4fJSXBIjMNRIravU9oSCu3EJSv3ci2wUCGcHRgLsutL6bT+
QwcJikLtmM5hIlSQVR7WJkkekkM0DvEvP9v+3YMshmV8z7sQbyI9AhOiozBrtjojrMQ1dW1+MH6t
ZF78rYZ0npTZcFmbRleRUWw6WsGh4USBZRda0h0yP+OFQ+4Hh0iRnzYW6JvhUj7MIpo2fZN4BXk/
WYxCNhbchUtA/3ZS/bIjJvK6qLi7RrAnfbGM0zTeTEM2QadFDVblNibv1MnR7y196UTll338MdnP
gy/aMUkr/sEGXWS6x3HFibdaO0xGCXKRj0jbC+yKEEBC9BYiICMZmGVoWYMeFCw4Ea0KiNjBdw4D
oEaPuR5j3M6sbaR481DAtVofPoqP/aXlfbpqh2pd/i4gIe/uw7fGBfwa5NXFugFiidr3RGfY5f+9
jgRD31f9NwSQjAq0xclxXPrpWD7gqU7B+3YiqD6Crnmm+owm/F44P+gl5i9yBybaxHVI17NFdBEk
kCt9YHTqL1x4yEu0TiGPguWs+YeyUllJZbLFFqF1s7uIPzWEJ+yPeUsoUT4KW3HNuKHNCDgRj/Ov
2zsmhZ6EG6UabWG1pbfSiDfX59JsFpTBWZVqSkaOPmrWabf6ZDNyAYe7bnvQetj9+gwx7p7f6ntW
jpgrB2XjYlrtKMGH7qOUAKAGjSjH50l7A2MHDgg9Uh8S+T2s1+uefSi+sj1r0g13SaN9epn4qAI7
FsPmYoJ05xA1I44rwV0flibOewQy96QAt4rqbQcSrWc/1wfEpGyJsB+sVmZzOJzf9AQD/AmoGI/i
CwwbNGsfMdTkDqivJzPJS74abDOS32Kru2hHm3z507LoQjajp191xSQbjnewRm/OtZ2gfFrIsS2y
slFvnKBQKm3/oRhB4PabgClphv327qQeL7Meq/dvlJSJMa0rFjbL3nugvxr0m+uDl+Fm63IU7Swz
y97MtZroK0sx2Aywue0PQPqCHqv4JPXcJd+qUfIR8CVZtyVZ9OALSLAGnq1lcQlgqAbiQHGlUPZp
inZdVQJ+3nOq8ZciFeIPDEotnhfX5v2w5d8D0B5f9pW4dqw8/Zsi64H3OhTH58jNgPGDMXjY7CWr
Bt9f/eNAMEcVzbf6L0e6mdHnSfAUFSnhLAtCEIHAFYkP36hOHpFF+YM0utpQC4D5wFQMJm5jG0Dj
earF+dmgCDkBvjNVfW9ZhjafK9JjwcUvspYbX56dqD4eIPxhCswJwS3cmpZXkL6hKkmv0f56xVmZ
7PIbsqgjRDhvWJyTvRiUK5VvVETr0QUy2ZWcN+HrCYvQF4SXlGOJcc8NwxJ1ZIefXqRCSA1LGaFm
e+iGYL0nrxXaOdgVAQ2AGKjwgxapBCFZ3AZI9vypmZy+OU2343v0wujPXUYEXqEeh6Dmu7iNN5JN
o+KhMtqPZdKtYZY8R3nRw7c4oO9S8kQgnJXXikQIB5HQxmeNqaNwJbPVOyKARTW4n5fbdp1vbQjA
UYcx8sBTvtvFa1q857bMDwKOdI0B7xnqAo9wkdDASe8YXRlRRCa/lYEhMbbO/Gp4SxSa/0Rh/f/8
Rw+82PUCH59CPhmhiRZXz2r27jDJ3lKC0RjJAjsjIO6oxf5LDIqkmAlqvzQtdPMzbU7KIFyoqh2D
RO2hTKPAZAtbi3H/3W1EPj9wUADN0YRoJSc8+8Cx7A8h9f7j0lxTlPFaTiC6xS8rZvURsX+p34v6
NV3FaP/kQbTJg0khaJ4OSXv3hznO3T3UzYxrnbtrNLPVz/ApIJwh+F05KS1Lwfm8YsGmTUZQWNuB
phu1NtYBHj37TrS+WBGSIXR2T5Z5FREkC/R5bvMQmtEtgkcNjioXHN2pddq1mtpIt0SQig2S8Ufl
TpxwXkce3WK871fImXyguSobBLuslgSMeZnEm4rj8o6WYPdKyr5JjpJseVUjngdxFFQHnxAFCFAc
oGmzmI2i7TxMQlgBGQuk9s8KcObZuRUmRMKAkQ+qYekNPJMiOLK2u1BTty0tI/I+ZLOWfUKbrdBE
5Cc2uSKWaazckHWfQ1vxiYt6VRbSdhwUXqpeg5W6fkUsFrJMWAZZSRTt+ncLL6RP4G0fK6IXPE3q
NWPLoVCkvVOXMWXhJ0BM9JpGGhK8xeMV3qUZng13z/h3Oyu025IXwLVfEpr2T0hdJj5qvNAVkmcz
GQRIHvsbrntW2h95oXMTol6t+naILT2HpneYchzakHEC720JefZ0S3grmA883xWCDdNvgeFlI0FQ
Mgaj1RYr06K0cNM+UhJtWAQku9J0CtVNibXwYwMP7qS8cqpfzlObtGZeHRAU6Ma5DzT5aVfC9hfX
LJme53h3qv9/5tgEZVfqcknZPAfb9htJDKIzGW6zy55rUCYZRfb6QvY8ktYNAJp0jJ1OJTMyM2Ia
nJF5+6VwVuTNvAVC1SWng3qftE8etiKhmZ+Nh2VPlZxKJt4WrbROVAt7dq+lPivxe3ZfSQ9lwqpW
0SmZWsG9t52ZhmZzlK80vEyDAwOXEm0wUyJHXcFz4CFhM5UYIg87g+qjWBFRKxbxki61WsRMA/Fo
HGDVTYD8iSldDhZ4VqonY4vp66xu4fT44ZOSDMAIlrH/C37nW9KVxlKSoHaMFhvZfvVzuV9La06l
u+W0LOxi/+J6ve+KcyomtlS0XLRw7uNXC/ETlnpt77Y7BFUS75LIOUrNxDcM/csGG55oDkEeID/1
myVKKM7M5Do/dB9GiyqMEFbkHbbcjzRbpFGcGhg1tY6qF9gtivh5ZcHzbkKI54PWETeULoXPCIzK
zw15EdVqfrCxayut9WMUgtM3X8Rshr9G6SeXh08nnLg29UB0BvUm9SB+0vB0VmIm2FTgRth4BRWS
IL0/UffLIt21pBtbK71JiBtjMeP32JNsFTKakoh5YvB9wAnpvHU4hpYz9JHcFTmohJ3UYVxBSy1R
upVpU/8SNkv8CAVo1aBTGAi040bo5YBZ0fdOPhcNFoDPczUDWiabZdlbBd1Jop5rzrqGQlK7ZUu6
5yxEfozMiYeySmEAmhQH7fabYSENyJUAX9EXQXN3D44WP6WYtuWL/RphvOJV6BB1ARNlQVBHTz9p
/rYRxxKvxo47teguHEl5mP4+midac+L5lvBBbTNhhYgBmQDKbDKo2etT/paSLVl0bmVfGKbAMkIG
nEBMdjT5AniXnW2eQS+o/s6cD6raB2vYSF/aT6WOeDhSFZAcHIrzGTI9QWCwMYOUxcrQmZFo6U+U
4M2EyTkQInEooem+dTEWsh2U2PUH4xtZZlPapx12ithcAtnX8i4oNaIcrJbepvLOvcFvZIdxVifM
z5kNl/1mEyZ1Z3IMqXLVmQfgsfzznBYTdncqpaUJop0Sp5bSinYtDUBefLt78RhQMwMq3JJVuguY
a8rtHee5jvwZWuohGG0Qj1A79XAh22TSfBbYSjXSsSzlqa6rWT4dwKOzodeLjjzxH8n1P1l/6jYe
fR1jlQiRCSxPxnR/rqHGcw8ZYspGlWZeuR5L2KELtUBF8+Jz3b3WGOEMVf8BKf+7R3IkUZYnYGIg
7jy8AQdW7VkSIBppUGekpdXzjR5kQnSWnh/ufDhspbvEamIT9u/XNJwprc2Kd1J2mulUO/1b6BlH
M9IGoBrGDfZSF6visJtN7Mz6FYnBkH8WouRybCLEqBqMsvvhJ1+N3oTCkUVnnCfJWlnG1fbuBrH/
5E+xiERJjdh7Vmguakub6Byi7KOpntq6GbieOl7zW7P1k5PFxtNRoMh7MBFBisJceWJnycmrA2/k
bhuFTXBOxHB1k/KId3dcpo/l/RwGDiwzponNaQACN+XzBgPrXzB+o4Xumunr1FuOcfSZJnVfUf/O
4iigdGHxRPytmmljfrHyb3JlClW6+4/Q+CVVSrMBAG3B0ql5Y7NbstXmydXg4HFNND/LsRE8OBfF
ZP425RnsKiV6MMPUCtZP733/UvwibvhllF0bhS0QOyFrQMncuf8GIsRxfG7q5tah7Ldh9Y8OFTyw
xHFm83Quq2jmxMrTuUY0dUqq7Fi1obi4mUkbtKjI1RpWQNZmjNmEUwj53/Yc9OZiDmCwmcdcHlgX
55isE6VKsHVCXUS3dWzrrqUtQWTO1budcE0o8N4orsn7yKoulJIQUF9dw6OjG+931No4QrCe/P5t
AHPHT9tPtZ23Bp8Gvtf+7ygMRapFF64a3swBoZ8j8jHYPDX31D9ygCgyX6k/ZRvtERJ3clgNvX36
4degELqoqXy/7tLxPDy4nb0XwJDT7H570pZf9cuMsN09Cu3dDBkhqysSf8vnQKIs57mRp1r/fHBE
CuK2f13SaTje5BQym+mIZfesp6rQAmCxqMmkckTo5C6ehfjvxCStPkMO2nIRtdBXOXKE+JUARFzD
HNA4AAMah8fXgq1wzkB/o/0xg9CfIrERAn/RFBCP5SSLRoVuZ6iGbso23hJvdPzgjU3/0eNwNpWn
PpBbDTKbqaLLpgRwNMyWghM7R6sDaiupQo2JOxfkr1Izy0xGzJ6017r3jDtZDCjcOJIcsxgQCdE0
kYbtr/8YUS593k1QONxhnLT29g5O+QPVhIUvdbzdgYm39jLuqBnSYjQBDvDoxWfXx5My2CrSaVZi
YlxrGr6q+jHBEDTPXaY1ddUe9LRi/Fddm59rXAvNBetvZL9biYysUSE5KGzpdrmOT5PHpJuTEGs8
GmuxIdKiviS78WbVoYZ/DFfAFq/JB1QFUPspaB5aNHvNeypuXzCFRH6KugqWDoTpYW530b4+qXyf
f5LZsKx7wLt+FmNJ28QKUvz75CHNTuPuzWsBQ2P6wRQgYhqPnoLSXTBpEFwGSaiS59CexlKaslJa
KYyQkavhqwWeDy1O5dQUabnOOqb1ZwqStkc/3TzZdwRIq6KegvuQpB6Dyhx02/ggwD4VF+cVkP8i
OvgVusRR7qypYP0O1uQB9W1Ek12ZjpJeQq2g+3uyxIdf/3snyk+aOnDPhGv8OKslpoIoYzds089o
mTNMkMjEEVBJlgGy8AylYYkxDeJ8y3UyhRAlhSNzlf7fPGW5YdWQqoRDhCNDQ5rklVTffNKGM+EZ
ESA7ZqBO0yM4Q/u75Zh+qLLfH+SP+NItGfx0BelWc78E992EfPGQpUonzPK2eV5Wqt9NDIndFppE
+zoK+SkWhMSh+bTIHHjyeQ/k9wglDKoZ/UTvAjjKlQYPX6G292N7qwy0WwvCIPXNIpr6DiJThHBK
WUiFWSmz0chsmq4LLBvCk+bW3mKnImtzatluNPGXwEZUZgHpT+N1LLEus+aWIFMR2oB1APkcMO92
M7fLHSTQplvsx4iPeyjnJaW0vdOpsVJpVbFzdB1i358fojo3+bgMU8gucIz0AgVVYEHYpMjaDNgg
dpuBmlicZpJk4MN8cLnkakgfh0R9WDjTakmcN6SvUgvuzjpI5eKCSnvEzODOXghpMjqOwFYrYgK/
kQhjy6dLkhyxQwtUEqdpNtwhqlYxzkBe8hh0lipAzQwor9n62XWz3gLErtUHO1rQd/Y/uUVYoyGF
XSDwKx3Z/Xw6PROe3daaNWorhCp2+tFQsypC4Tvd7VQOTAszc5b+D718BmiJsjasK3+5QvlYTPgY
Q/UxMRgD+a8bwNaBVRQW6YtZYe1jk8UsBJxwMZf5WXPY6s6ahOzG0gZBrMLIiWSHydLSm1vZBx1t
2+tkTJsG7YuqZf/uD795LNx7oCmNjbaf1ZuE+zorhXaH9su+VKYM/QsmgtR4FOsMHGX1GtiuUhZ7
pUyWs8RS55FpNfn+dofE2ywAjGACwk8Ec/a33cdZ89Gjd33WwwZDyBm0kYqTaXTTl2wwY5CHYnNs
wdyNrHVioF+WBLx1N4Oh84bzedHzR10ihdfeXtI30GZgIcrJhfPYFth+UbgeHSMuxKJh7ofh15t6
MpODIiVl+H6m+OH7+ZPNqeJhrlL4/AtjaYIZnwGveI11NoI7Z9iLg5nXo0XWMnXQyjScujZc+1Il
OJdXgDfNAJzPHNI1AbMJJcmFjJo1ub3PjqQuR/7nq2KI+XuiiGqAvU4gEODFRRkSUwelYMBXcJC0
Em6qtWetg7Gvo8Z1PJGB/yNOYkaEEEDj4DADu9quSgLEPJSps6HZuE8bfMPZQ+ZwCVYRjv3LD+W1
tFAtYLV/z8HY6HPe7O7D2+hGF7pZCY7PsRejYnuHHXZj06EUY5qy2PgtBZB/xGyByYRdeEmvo8ws
FFWBY4P9cSHK+dwGVVNud9iwaEJN2dtVq+pDg8hbd80NvTO4JE8xKPaV26H0ibdEjEDg66F0koKm
qMweLgZNgqIomv2H+4lyfZvt3MGsLDt/ahPvmfks8Wkeu1O19UzvSyB5dTHYpQdIg02VML6GmvOB
eGF9LiAMns/DbiOKdv6JksmYsbnB1B4MNIxP6Uk1gLocQLmTHPSU/5gQRUvP6jqfXsC6H2V+yMAV
AiFOy6SeOU/QFJVH4dmFWXTuOd6LHe7HxhIMijmF3GaEL5an2aLRDe6GjBUVhVrKi3oJefXsGk3w
PJTW79GGuWOC7yBomdVLfxcA2WT4ru8qH1H7ZxXd4X8nbr1DnPlwmm0163YBN3MCF3eK3/RYgyxb
FRA8m+kUjod6jrIcu8VWJUfJ+uNMQSDA/tyWo80K7QpxsZxbMo58W6B/mIQMRgMizTuvcU0rnxKI
Bp1rfrhiYcgDWdbD6F/z70NPTJANpDj4is/SFARlx0boHS0A4UTyrvuNGQ0NgCKW4KekCfF+UZdo
bvjc3K0orGBjRVlvPfjCFtU+WV2SI3Mr3zBGCNgS4+lHI5ASRZBhwogSgxz+Y6mE2j3G4xe3epBC
2hNeQVqPAKKvihC76X6VuiDOenkNIPHogQ0de5jII0Of3FXa+7XS2tyV2Wg+6zHBADfUJiazMq6V
o/48LdK2Ap1mt+flakRKI2+K1sWyg3BN3Hhv4pip54fs75OvJVe2arGY57O0pH9eWsxcPDo1/1WY
sLGQb4mV1fj9wcQfwekXaQ6CHQAPjcNSGzPQxN56aUKN2D6d8iy+re38rM+m+NTAjpUHPwO8ziMg
zQ4I9Z7X2J3KpitzIpjxp9mX6uE6eaAmxThz+37D7hl1XZAbG+umRattQ3y03RwNApsRZ/2nCq3l
WwRzKnQFMpUtYvQa8NbFO1YQW9iAV6HOAoYWryoA0zq8x4KQ5vnpLE+TL+uS53yztdhgLUn/Xder
d6E9yAqMVg9A5Ga6oU79shnDZNYET6/ULOAQQnu+WuKJ8PSvdDheL/TPj8yhljaDogBDeEdzcnVY
UTG1aPrlWTWBVfRlJrdWNPudJDHXYs5btGqNo4/mV44DEDQ7XdAxK2M1IP9hiLnym8qn2Wlq9CDt
F5kx7ENS2BjaD2objZz5a74T39q5wC8XmqUYBs1YcesqGw/NdNVNJ9oXVIg5jICY0gHqu5I5IwNX
QDQsmdRUt2rH7G+ORWLC54MFKvA+/pEjZRYZkeZx4C7/jtjl+MNaHELuAOSND6O0w/wXNl5PjyhL
NHeFXgQE58pySPA7TNoq/kSSoyqon0EvEb+V387PUrA3ClY2TGMmyDsVKWz7cNSb8lCE92ZcrAyQ
ml8ZHFbzvVyHhfF9fIOturQUhDKtEQ3Q/4Ff7Dd2MH8iC7yqiGXP7q1F27SjAtPQqOUGf7rM7coi
fwjgEsicr/B0+rDmUs522lDZaiCcrwkVfGB1nR1zXaCu2g0KSSQ24jDmVVdHhJe671Cgmk1GwrWt
YbNOWrZYdKnK322j4/MOAtQdha22z9eccqFvnQTysfUmvbGEruygS0PmXd8pqPrVVQM28/KznapV
mQ6iCTaJj7SbVqpyrjJTzTiBq1usOFOe3yBpRmdysKRqkr1oCVIXB4OOdjLRwYJiRaMqOUbqPnoy
CqpOEJTDk64EP8WQYns2AWE5MbcYk4OXzG117FPFyu8KlxyLZ8kgUCObegrO3uhmPwzLsNbo3epL
G3GrC+s8nXRCLdsIfTLXgje0VNToy+y6GjgcyTutzHENdK0TBf8sfshv3qHKSkWj5o0QJJ+9pLr1
9IzQ1ALLGBLS8BkU1Vss+Ezc3ObG1AW4ZXitVfnXgse4VWKW4I3rFGWAWmiJ6XnZ71pgQyEcdrA3
v0Z9wT8Vx16kPL/aNei8nQ/+yIdYZ7OFVqHphfhXvGrGYDFpvxAyXEsHOlFw585uAq8aVEQvbnfr
2t5vf0yIYYj5UXfrvkdzxomwzSFS75ioFCq5008rg9zsPNFad6kGM1qsntkXnOLN3yTDgTlVvDX5
Ek7VfZyZorwSpnFOzIbDdgg2+2D/FZXaPmVfcrHVdTrNozI+rwLsijVmxW/MXnihlCbRBnmw50Rx
pTUFrtf0fPHepJIEd6Kx1XfBQ/kVfHMSXArlYLLDOoWpj6sNmR3sfimWlhr/5g5rnKC+9kgRfAeI
gaJcQANIh7f+qpA+hHw5jTBHc+zo5s4Qtp/zd6s0ZZGAwbK17dSUXZb84xFSXHtLKdshfnErRlIc
Ht7/GzFGuVBWGMFXvSGt5NpnzPUNrVEMFum9ow1iNxzSdp2TQoEumcGJOPYDHCHfvh4tk7dhWfoz
uNkkuGiWzD3qogGwgOmM+KeWFhFxOdCU3QYPN2mdY7Ug31/ko3EW9nTIAx5N3R1k0Sdtvxu6q9QU
o973dJV7Q1nPMe3PmP1AzrWygu8vp1Gw2iNea2loPb3oJ4yWXJNzKmIGycWpCBS/uJU+O9aC1KbH
e8O2GcFuz90PHy2k6PuPn15ohY2nDS8eRkoKI0dmDhXr7PA0nNwxVaRcD0MVEo8gpfEm3C0/DvVJ
f6Cc9S1jfcoJnk8WVcWdDeog0BNa35gJyqeRzUqpyQr5opw2vHh3gcRg+cUEltUUQC/A8ds6uCm+
bwKKJ0tVc98nXITqAivo7DVCD0l55F+jzBplEiQVaSFGAHqP1IwzrjRIL8vPC2KcqufRvVzBm2el
H60xv0T3x29C/SMo0dp9NRAvxlTQd/rEfw3Z10Mc4/Y2hBC9+vhLC1y/Y6T3dUKjN9//eWvZCU+/
tbcq/7ag+1F6YMsju9fp72AVI1Wz7UVDuJj7o4K87HAtz9vDv6L8a1Q4cxo3XTYly07Rc8dP4CbS
1LeBwmvvZD/hHjqi73NMoJyxcqLHGYOJoZIN9GRnPDpOOBaJhjqJacXbL17xsWR6FJOsemDO8cDF
Avp7RGerwNyiUswrURalkGGOyOiLOgrJQaOsoOcPuD/Zq4HWT4F5DnhIW1ZVn7t9x3xyisrqWL4j
en8/EmImVtVVIT/LFNurqWuFB8y0jg2ZZ56hbecrx8OhdSaXhStNXMSTnzKOUlZsDRb8lC1O++FB
fxHy1mOIMRbQf0IJYmG9OH4VxZ+GsA+dTRHUYlbnLgzJQuNJx+WMTCSxvGsiXvVkEGxgUokugWXf
qOPMIheignJZKAPfmdGu8qOqLdCoFn0zmQyHrbeAOcRKZlxd6CI6L3b1sIhQuxUZpQO4XPDP5MtK
ys75M9t+3ZBmtCj6cJ1bO8le9xq7itCXkvwXm/ZFpKHj7EIwRyJyrL2/dzWiaO/AlOiXSNSayws1
0K32M+TCoQ/utBaRiamH4qU1xT+asMe4fTW8PbbwpjyfM6Um0p5Lx/DFYRjE/+rTLVvUjXlHbeuP
XenPF8EUKSLWl3Lrkbepr7wxlr66b+yzLpW9TguuSfd8czVjGfGHnB7W484y8ZpLzqS5pKm+x3n/
xB0UsqnqtSiTcYR8Px6ku8z+ZDvLljkoWFgv9gJ3zYfeX2bVuxenFSyuQAFW9updQh00ld8Ovsxn
dsoJA6bGHYxQA9BGfwmnYpxpiCj4ZY3pw/acMOfQz6gdg+Y8mayZxjlJCj6zsQIqyuUB7N/EwxY7
h1tpljRieSvM6ejxgEYzOl/GcLP6ubuZuqO/PKYphDS7n5hATfJ42xgg9Vu0pTqfZZTHcqk5Nn8p
vW/CZ8xqZkSzHzTlxW3nXHjRfcs+5oiWd+0zh8SggFTuVoYxI3O9YF/Cnikda6d1b8QIbH2Zap25
IC1MX6mJo1N7Xs/EiyI/CMi11cwcVi9uIiZ6OH4bsNHxGCGkD9EQeo0xSu6UEuvqkFYRUfhuzGHY
TvABsjeFaXy7YvY7nyG8cE63HzdP9O5jcgmjxmPRxrbPBYhP2AKJcxVEv2tx7+HPp/KNXU4fy02h
QzIi6A+A/hfWtzxHc5984VQEoBky2skrBNVT2kBNFDBL5ID7i1iSNTj2w9JHi7SmD1h0h2lMNyhP
1QX14Q3M7092Vxhekn9RiAMAOXfvA5GyF8EC1S21pOL/ffEDkbreXj+ksIsATa3mw6KHs3dMqTiC
tpB7+hQGYvZ5EM4ab2YTAnR1OMqMpWEqTnZvRyKd9o66i6CBfMqcMU9sZRCT+AHjCmAoWETWBeI3
if7FeeDerg3ExZSSHu+WMM9qDZpRmaiZ10vLpaBZ6yZUGXgNBOI5gy/pDPwlnHbyhRh/gqyBlqXP
AN7yhcmKhe6fs7sgTxAz0dtT5dnPoRvE1NP4gjZJtiA5cjUNyoLzrgx0rphKCM/ogpe7Q87yqfZ8
JtI1Nd5yfrhwSBmk3LNKgfhkEmDQRtLyM/mU47WVCH73mKInJJWPnI7JCIgXtc07DGS3eZFwJEWs
8BPkJRvfBG6mAcSH4YjErc/HNkou4X92uAhI3Z3qis6QMqJoS4dkXkfBJ9PUfCm2ZKwE341d49UX
VF/aQKG/Gwi/rW/zrJv3pKAWVOxE04UaldLyuej3kXEKtLAR3HTsDFK3eS6l3RyUcMLfAB8L7uKk
GT5f++ZVwtibKCRB98VcoI+uWmrhg6q1obx+BVee5a1kvTHMf1BuTvYM7b39CVG+PtE5L/5gW8/i
AqWl56SqvpS5Whjsz9BX+0JTmOt1g0Iovdx7iiGHlZvtxTsYuc6k1j87dSm3qenq+w4huJV8cHJc
Kw2zpiEXa67QfZN0QRRO0tKKcEioRbnQ98j8lweyjs9HZXX12jrCfAT7SQCBldqON46N02susAg2
N+o1z0/h4Zpue/QQ89PO3PygGxO7q1ngRo77XQMNNMQINsu5HhQouTAhLgzWv27CXta9nK+q2T31
dA/Ue+jbIFPVA1Ue76dEev8Pjd7dXgzZUQ9dYScsQI+sc1fLVpqr6ygg1zubXkINpUxL8Y+7Oll4
FDD4+W5/zfY6xdSleZAkEgcmntOjSWKGjwQcn0nHTxTf8LSVxWAwa2Nz9HbBYhY78i8NvhLjMMp5
fMTSlze+BBX2dqAUvTUvPdzhtbneOaJyqbFWMpwnimlZY+Np+7yKmHEyhpIJuxS+tnBM5xW+LXjq
Nmdwlte8YCICvj6o6l3nchTf1Sc2cbwh5bZNkL4cDni/uoHtEH3Uj2BYaZu9SYxyWK96or6JlQED
yW3I171fYspZNYMBh4DkBao5SWv8J5cd0BzWEnnMymUg31AMD0/mBPxOy0a9fj7a2YTPE6/HfJoB
TEnFadNhCwEtyy3a1OLoj8xIWLB1fsMkNSYoK25AwXIZrVbS2OB4Uo4FL8D+7dyQGnaiaJd8dIT3
yil/0Doi3SFbhsj/lioxr/wqsUPCGqUTLSSE2tMyiqGQMYrIcBm91SaRHZvz2XFEGE8v0zzRwh+y
NT9BQDf43+ZIt0KtU73TxRTmmsGjnp6tS13na8bCY4baMealdxWhUOzswuL2HpkIsTQdOA/qrt9w
asEsXzSMUDtJzTaQCUs8dimtjq1DZjonx0llmqkfig7lUHt4THRIl2/9476Gsvxz/26HYkKlaXFn
4963AdQdjdtRrBjVzvJm2q9dcFnoV9ou2nadGY79y3Rwi8ONvsWes7D/RUDK528OOCcWD/tcAdL3
Wdbv3GyghaWFeBS8cnWyHWlqSkvGStXFj7d357hpuLThzzUGL7ZX7ElahAF+d9HhqHWcygQfaUFO
7t3e8iLrvZAu26hjddc66lLMOi1K5u4SkRMs0BQY6ea3l3RkwRT/oY4UiqLg6LYRU9XGXG9MvHXn
oi89FSLDhN1VRwxAZ/nLTMjOEyPQLKUXjEovI06UqkwIXYy+HX/ykAoMssgb/16pOZPaIhXqn6wq
epR4lB5oykIwfiUmUXlbmoV/r8LQ94XTyqn5JjytKORbgEaJXiURw8BvqAm5OwlPVP9hQg1gTpqy
4sMVEc47b2UmgKZhjeBxXlBPnGXmRZgalA/n/SS6FtB6Q+yCyUZKtF9axYDGW//8P3JUqHV/PbjD
qnNbFGDrEjwOx9lhRW7CMdSjhM4POUE8SCbr361lIXR5SCThrh2XpXXE1GchW8BTtcqBK5FG4PJB
58j3NO03GSgGUzGeKMy+xnrrob+o4BDtbup0DGMDowIMzTV9FTUy3zxPXshYedXQmpVXU+zpU/BA
SOD3caw22vTys3/Kf1r1kOfM9fCI/HEyxIG94UQb6N4SDG/BLWdfBZL19p75hMco0nXC/Hlk+Z15
aDiaeksJPazjWJYRIhpI4BeqjQTAYrvbXXpbLogpXZ/2EZQnrhNS9gJ6dlBbLF7F4jemyDID4piC
ubRgcCXIIO66t7Uz/hd6tgsIgB+iZww7zu9yxvIK8OhkSbfmUgjvtaMRb9C4w7mYsy7N121yUSEF
e3Bohi/gBnU9isC3V7e+oncYDXWv+3zeoDc6JrKxUzYaTBWxVPS7x4+h88GlM4oons2+znhdvaXj
qnjDvVFa1f2qo+nmChF7+3N2L75d6LoP7hkhELxnBLNPU8eAewzmlQnE1EUPrZG1Z8SVQBU+Zw51
F6VsEuf2tgVwenaTRctCt0CtTiLJyO9U203DuqkkD+AFpfKjNfzMR0fxmTfNsGJdw9VtLV5XW0oR
2f7+2rAO0CpTJ6yQbSWAIeqvgaV8g0T/b2xoyiY9B95k4TgH7rJ00W20HcFqW7XDYIJMWDMvVPLV
PaasUSZ1vmT2IKI32rJ6h9lnOdmf4oeWQwBhihMk+tkjX2o/g8lrH8n0X5mTwAPG+0PGzfHjlFpL
Kx69hgCQmNOzpWiIcdW6jNRXx/iY0NXpnxBTdsJILxOkfGYIoMPLdDMVhlIcqJaXP3b67LN2UKMb
vnBlS09PjgyZLj2X4gh7mjj2bgod0oAB1lsJQj3gv71aFZIvECbQWo+2puyaQsRcT2/S0CuFwKAC
hAuKn3y+BJ8S3gQ6OIQtNw0YpLRrezOmhZJMe5qlkInXWew5b2gULteQjMjutfTBn4BLi+JNnPnx
ZlgQSn0GLExt95583G4BFMIG9+jeNCi8ywQQ2SY8t+/Ysx+sXRIjgYSpLHIHSnr9vQDeIqwBZiHv
XdIOWQa/dcvamAeXJs3WpQkr51a+2uezocJsLQmOcvehWoIfLjZIjF/G4d9KQnr5gx0bhSLK92CL
gksY2Kh+c9kebBP289vlOFiHYyrh80TqNdZ+k5XmDG4NEkNJpWnqq4/pZhJhjt8ifi7MFECejc/B
i9L7vltN7Kx2KVYuwOV6rjlUvT8C6YefgD9yqtEDxUaUcy8G4jVPGY6f8wudV5USGLAHyM8pITpt
LehWD8WoyOr4/4aG1lovQuNhPHPE7HRFf6kz/IVQgDf380ZX4OojXV35CqW8TRinmNm9Ax49jcBQ
+GJ/mW+d0VUvlSXfD18FPLSoycuF6+HpCImW2NE1cbYyN1F6iAjunSwyL9RuMK6W1KMH+7WFcwET
yBQfQioSICw59++wdl69/9PMuzqDrN2a+nTmRputrsZA6XCruQSYpbm+vKhDzlLJs9V/aeT1SG0U
NKriCy6rXp4zxKztUvW8f8wrZ0+k9VySE9BCkTaFTeAUfiSK4mERPSxIh2dB3Soy5tjzx5uz/Sal
o0Ol3+wU3WbbkgNQEasVimoc/rgmhDTIghMnW8e8zczxopl+UyWoX/og8l6diAncfT/xBvO4Psv5
kMj7MZ7R2q/0uNVaBUGNh7ko1LwsxoOdbpi2ILml4xFMlCTfB0SB7NPv9z0gEDj2X12XPFAUuJAV
0RD0APXZJD+8Pprv98UWtOTVVxLW00KWmHbtvftArIqoAShWhKrzWMfESIqyKueWBKuX7jU0GofV
oIjAo2D5nqu/cK7tJUYSnU3BjAXJOBSH7zF/TYSSixBrHwU+D2NHPEfpajKy0nfP7iMi5iKZVZHx
+bS1QOLx+IkweGZ0OCjykCABFICG/ZtCw8u8OqameMvn34Nr80sqTsK/4opgMnp3w0fDPNx6gsN7
jJFmG6pb2jtdtpWkmIWdWWVNhAxEhsohbsid0zizXmYPJ9myBxxzXpVNMjQfyqdejop9zG3tGdkD
VaZFiZnC8r0zFVUJRfLmHDWTCgRMQVrn8ozlBiI+SCVOT9ANHakynmoMJ1gSCwl6g4E+IH5JudCR
wKjhNZAztTczs3pQZlzePPPnaIY+lz8BJuWlN8+fhtJkRTlMnZcnzrS5KNgW2Iuhok9QXDJr4TsP
7m6hp6zWzSm2w+LIjOotrNkAwdtg1pLw1pZkGpNamrw0pYvkzSbZbIi6Ih2bfq21T1gO/yaiFs7C
DMgb11pY51rehO0DOnrgppBbr3aqBWDOtjvsVQBsvP8vReEQ3vVQLqkARfbmN8hCFscpleLqIJAy
EilyD93J11JtvHuntqWOQLQeFfa7glqZ6ly9pZv93hsBR3K0Fc7wVxiXBxq5/yuqYht3cVM6FnwC
AvUaqbKcbnvmfSZkGYKw2Lp8Qs9MEici3O7vNY6w8WufOCOQm+odrXUg3N6jafg6SwmQZOLlj4Bj
2FdDAjjZnwnzzd5GN1ZaT1hDu3VZXc64wtlc5g+59MjblkCDBIvn1BWkpQo4tueMltOM1utvukVU
j/Kgowjbv71X3CRZ8c7IxnTl8lvMsiZgDiD+c8Im8KSDw36NeQ+4JtRnhbo03Bp6S8HOK8+eP6uG
3StezAjORYzXW3fIcSMPkwW1oxV6/qvaGJhHJNFGqDDYWK10G00wj67Y7o8WbEyVcuvdzL0i/4vp
tI8xLGIvpapTzSFHoiMXWbj3ft6OvqyAsB30gds0jPJLTT2wGiYGr7sUuzLZwerGoVGc3zh0eDSn
U5pfgatXSWiUYwtqKAK0oBPh4Ncedgxodpk0kPWVJ2YCczs3m2ZzvgL2SF4Vi/wy17eR8zOs7Rxu
rnyxsye6juxh0bWnZrIlN39n8DZK6p7CMdT2tYfHptAMigICybCdFLQkxe0z5Ms4s7ZQDFWy3W/l
PzXtFuDQl82kBqKEy20P1G8Nac8WOouHUxEOl73mt/hVNY2NubJMwK74eJlBtTif3RTh4BuvdcHf
M6J1vElKhO89IeCRr114I4c+lA6lLP5U5Z4g3cDNYFfAG7ClqvgKyij6PSu2ABuoEnhjbhM8+XDX
QV2XGR23BNMLp1BCm9sCwzvvplyuiTGpu5P1F//t4W+CoaQhypWyU46L3wSDc7FjGEKkGP5pdkwH
9s750Co/xStJlreb+Sw2kQ2ERHhNluwSpLY6RXYrDMHngHagEEylqrPg6ZDwcGT1mpiuZ/etFSnD
sEoVlUyRGRgmnpTNlKGeCbw3Q+Vi5TEreWRShKwX9zXCZwpmjcGX0HT5AJeQolyqmDs+m6VOoxiK
zrCJGD5DBbgGxm1UYE32BTtFRVeHwOPhfi2KfxfGYTgIJbt1hw+5y5BWUeizdve9OvKvq11Y+q56
3QelOrn+kwj2HWBTvYTjQC1HEVSvIbLLXF02haF/wzvcnbWRbFyEjFcal97lLfvK+7/1qc/kL4t5
+xNh1Wf3ta6O6jaQNZh0O7hLdrZODNc9rtQVwP+yDzzE/MFBYntuZM2Xkjtys80J7OniLwekJIMt
XrB5NdtlCRZU7A+zzHWf455NtteVZAsELJdqtjJrps3rdnqwGVHnBXpnfzE0eOAmh2shsM0FyXpT
qXSO8IvQ8GHNZPxVQbtKy6aPPXOmIufkd3T87SC7GdBeAqJhCyZR2IkUf+e090zna3yqA44y5PMq
ui5/5i8lnGi14kiCjoSA4s0AN9m+cNH78R6Cvk0N6LJ8WtRAGATXMRVu5A4TMPmPeJWx/L58olDv
AhB5h1SJAlulStqL+TFk/qDx/yRwOCUomyoXRNYnaP4qsdhJd4FDkArJd0zyPkVr3ctgpqeyQjgO
7RtraktqeTTcQvcbaDPbWRGw0B6n94iYgGCpA8zJKv++qgnvgtAS1WyJIOo/rkhuoAUndRY5g1v/
+1ZLxelCW3jCtUvY5ca0/9AmAdtVisVQfx1q9Ce7uqWPD8jnv2PVIslO9SOMZXIS6YRBtu0+s/JQ
tsJMLH1emVGCE4mR5BqOkHZYmhhhTFtV8Sig/DvGjENfG3h7KNW+47S/YuXFHBlEtYWte2hf1sCH
/bK3JwQ9mD4MSLqJ+KXENqwq9D+pGTsPL/w4ihXkh1px7prwlEH+UHDOtetjcZcmsh63vzYv+Lvi
+zBZo6gnyFPa6oq1c8zJZMqfUqtaueq1KtbbYg7CALHZ7hx789GlHczLXtPNMNvrDZ0tcpr4xQ21
azlt9daAGsR+OYiQHPkMhE90zxKRFSDx+dSOyuYFIactptUZuyyWDRliJEPNjtE8n+V0NGeGFkwx
CBANkjXa/F47vBqS74mcPmGGfQsKVeXrYx4XqCs2mzomQskKx8u7K/P+WcpguLDsVbbxAHUfNzF7
QKryRVIhp/eAcw6FUqCERfy6+fjODfkRMvuzJeEpUTM/7q/kebOarvdFLY46hwiO762wKISVrduc
ChzYKLSKuW0Hu5kPUxL8BmgOk6aB+iqPWKkJF2Z+isbucEUuNNHA6MiQgTwpTiBHL2sJ3dG53jXq
s+YbwGe8ePU9dwXELb4n5ZNQKr3S3gec8d03moLqxlO23Bs4ixahDwRUqJWqt7k2A2AkwxJqXpB0
z8a2tE4MdaLxyUjdhzfIbco6Loj/EKB34RtJgdLShX3BPxl2P7D3qfIf0itoXOg0abaDZnkpZRhe
/iAHX1Hw7BVlTCG7CQYAI3bfexfPwh2Z0H/SdUGDGht9ydRgi/necQ8jxa1Hk0X2onvryObkU6UM
jdV7vBYKwU5aElR5FTahSdqKUCkrcS4YLlX1tG/TlNqFM35wAHWze3yULPecI0LPzAxWCXMW630h
PdV+aPYSXbGt4MvabPOwQON8AfrZvQU/fA0RtdatsOE556OQ0nbzFVFgcaYs2RGjTXqRNP/v2amy
50pygpOGL8Wyph571xIe9WotIalCHqFU40kiqvlANO3zNOwo7bPv5yv4u3xRhrCLGEdrUtgFv5SB
Md+L/Dr9Aqc/MD998qSyrPtlXDonYxYti1Exl4B8XfQAup0e1WeYoMqUrTngBisUa1WJVplEIJT2
quozuzIQszsIQdlRkTpfJbKT8Lh6Ko+Y+Pu+ezDdygRgiIQjc4nFcn+N7J1O/hUsrLDavedvmco3
SrY6FuEio0Q6/+2L9+PcM16jlrWi3u4FgaXE6sA84it+Wn/cWGj6Okb1NrFygibJB2AKp610tVdG
ZyrJioQn1/yXrNDtkvjpysBKcadmEq7ZMkThZXcc3nPtrd3WLw5xmjF54kCQxQjTOWmxqziuqXbW
iOE+m/tJ3hL+s7e3ngNNZ3gVYi76/EN+7HsjFdxBRq6ugeAI/sJfxqF1FnQPDzLhQFqFKJpb/tRT
XhO8Rp1K4g74xX3omlmojkCOYC7FmJfZ5yVF7EUKNKMeqjV67lpwWs47x/vAyAL/Ps6hguhEc5N4
dj27JndGUUgWRrg5E5uPCSOgYytPJmZxi+9Z9EGXYubgwAHkCgkmpKo07A6F+/zNkOxOb5dwcV0U
8GbD05C3EsqI+NXO85tKpNN/AsOrePT1z9CmJTvPS0qWWHzJOL4CmISfwurbs18CPN+YUWRHzbBX
pv+nWZAYs/LHfe6pRW4QnfLzzeBUbHHA5BX+ac6b9P3W54HXXLLF0lWzXT6j5b8oMY2Tjws98bMV
sBfbKT/3fFrOhZnRATvvshz06T8Txqcd1M0Be7GmRJegnSK0sZLDdY8WTEDnwdIjAgXNh/PZQo9v
6pH3KJsPd4zTxjz/+TjT7W4l4Vw1a8oLvrmhPqsAC5fcVRTvGNeBbZB25gph50mZ6E/aIltGfKLq
1qxQw37S0a2S45xt2X9XpWjgLG5bBqyuxkaL9vCADjF5uuetVcRZXdBSqBG+5/0HYEtSAfeFW4DR
lnc6PFK6LS1DQjPmAyWwUT+JNc0CrSl2RzRMczC9vGLJmjiSS+hBOccF/S4qwsIS6P0fjzBHnIV1
tS7X5LlpI3Ky5voSvG6p0DdBOGLZnAVmVvqDlRcGgA+okxHjzUdnYieJk7j8X0MIZSgQ4b4Maxmz
H0rlZiA91e+u3ngY2CZ5R0whjH7Mu+jiFnH8N/24qo1dspS6IXygsbVFigFLXrXeYtbs3qwmlyrt
KdRMdJF55w4+XtXjrjkHJaDEGYUHcI+XXQkMTdG0Xj97YvdPpXXEdnijuvGvX/4O890aU0hGDmzv
P6Lbdgh4Y7QQJEJn7SdbX4G35fi0iAj+neTZeaB3ZV6W0LjvVgOMrRSzeZwUM0ylsAXIo8KZ4qC1
VTdV3GAzfebbPYbxiwRVSnQZN55S7UZx6MGLleNB/rWUIHcrw5xiJ5TEM++6eGTQR2e3YJxyKAIu
AdDbRYWy0v1jnFg5iQfaC1DRPuP+bOHFkurME0rjkcYm7BwUL3BdhWps14o8jnpWf4WdX/tTSZYO
7u3miYqEIke7tiDE7PBoD8Q+xvAEQ0wLacsIjJscZV7apS1JNXkxPLndfNOpSahyWWan3rQxQbqg
s4kqOmGGMv1H8pUGLgX0MdHhcU0Am8xeGVFR3qp/tsL/4ukjC1Epka5ip4gXVzsbhgJ4QeVgKagz
tIiK85xAOgWiJse5qinNqqwIuKINXaVdIrCyWymvCX3S+nZCs9oC5lS/WIsg8RvtXHXLkmgjhma0
xuGfL3iKqiimv5F/t+Tg5BP4748bA41j2D563xOZrlTYvVVdBRtgmvqEwTpKtL7T+gc363zlJlXN
+QlwMulcuAkmHzIf7QrNKkcy6tqKMuiF2Ows9/lXVkZMXANX8E82qMqwoESgvL+iwnho2onzPq4l
DIcUoMNYkWq+zv809RBt1HdX5O7jJQlfeUMKlDKHjk++1ee6hZpY/SUZgA34uqL4z2zZAqMmn9bb
ew3MryYdS26FdbR6mvgO36vdrRpzs6LCSFYwJAFZgCDkDWjg+dYtAPWMAT1nzF4Bd7rdY68nEikW
oO2ryCYwAHqAmWlWZOJz8qOFVszkwkHF7CPz4SMppxt55QH8FyERZoiL8lzFFhJcuC3oQP27Ywmg
c7O0YsWzhwhum0pqoqFY8TjwWQ/czILefHcGx2qmPS05S/ItU4FXmZ17/5fFXrLcB65HcMmgUtTs
yUv5dCOEaue65Hvtav6KtsG2PKTUKT2LSyun2sB9z15Ml90PC2iXtVBp+F4EJ85b2rAR2fCjHsOh
AyemXlE5WZJT3SVJ3I9+VBc3pp8pUQYO9SHgeA8RrhmMqor/ZaNjgM+MHYNKvGqoo7z/Z1HfM8ko
b4MF7LgWwnJJSWyjTyxghACwef2czpDnFG0vqmliASKUv2oMRd6QDvcUvDq+0pzHGXBCJlvOztN2
Exst4bM2UlcnS/E7S2v3xl7xHAM2W7E15jZOcoJ+Y17UYZqguo+URSDkF50Ve17mcJpoXM4Vl2FF
CwtdvPu+u2Qbz75jRqI82h9y/vorU/PFwspnE9pW4DH0iDobUPoL5cXdd73pKaUNwH4WGwILnr+9
BA3gEG7/C+ahZkHkXG5427ErYx5OGDXUrF59W2vuKi+7DfxLVrnmJImqPgOjKIoyj4HRY/ODw6Bm
EOWcV13mtTyDiJ7S9Ny64veNIvihyG2PvHi70e+Rh96lt8iR4L/bsXgz75EIKoZMfwr6IdV1Dndx
DLHZHdgkrUoYXFJlAMyFgHX+ea2MBVs49o7vXtsb6JQO9wkmdDzy4RTwQNp0ActUsa0hX5DhrHqy
XAKwZbbNkriyX8dHWJEycLS5JdZsBxufQDCWQNIIOmedws9MekyuEGmZYrtYrMH305YzznIZWwE8
6IeF3mgA0uDLDPneZxRo5V4XJLT/kmU+PrX3q8uyfLFj+XFL/ly8avDIpCVNS6SFLgLS+5OaxCJS
ZEkx8W0BVIChr00gi8hgFFxz0JBMLwFfV+7HofqMPVyF5BeGkGX/wCLe1lPj5MGpdEkVZh5ipsUw
zbz7sr5DnLDCk+D0049KGgIcJZYUOVrQDTJwS2zsTRGJIsVjDP8bjlaPCUpYjziTpL53vEL5PdGL
VvA3o9RjeuCw3iWdHpjvs8fZO0+bNUNaRHb3u6sLN4kmpKfzzksleXT9oXfHRk6U6mBSeZJo8nBQ
ubaQLRxJxyEVsUrivAesFch+vHQE0kcDiR6o4pG7xJX9u1ZTOc9ZObzXAAU4QBuPHrMV9ACZB3xT
n7v2t6U54L1LLNuCoUInazC1MghYjvYGvzON28MHCkcDKqzLJwBn+d3vsQqA5ulPveZsvvgmIdB+
4F0ss7JvQiJdCS/kSys3ujzswcUZU0t/pUDwjTiE+n5GMC5brOLl7LEARUPpEzAZYlAYmdRk5kA5
oaf+l++woSMxJA6d21tnkNeT6jM/vrr3jBnij2dMhwP8Mqzu3eb4Xcjnood1lpSjrrrzu/qowHw/
7vcbtpbfwQj5pA9/WOQlgBUxwqQhDOqqCxmYXrH3Ok4bkEdZ9xmnhjmq9CSiSB+qcInO4hHWlQia
pNKyTrLXCx7Dx1BPbYDBjsONYXAPYJ5LfFsx0xxeG8PW8JQ4W2D+FxeOORGdhHFZkCQqjAOz6DOU
7+U78WSY3XK7ZWo1lp1oj0j0Pndo+5ExRgOv0yjGDGyBpeSLzIXx0L34okU1zH4ZT2BTQ1d0y0bW
gJpW+BDd1OAz060aCzN8VFgdjtpYPlGOLjPBByTg9sZSMO7h8vxvyxPyBgisQUNJO/Ouvl6Qvn8l
cWXmIbe2OTGKO6G/iPVyBKhxa5Bi5TncrzFOZKjy0ZouIkkYgH0FW2WI04KAaIY10zofdb/ejFHd
7dviS85bV8byW0niYSjSThBW+8tA9Qy6Fy2i0rCcdVcgG+psTEqRU3qXP+rPMAOJf0E6n0jM3st/
S+pX0irif5zCJtNYsOmMnUb6aal8u2H9JpclAivaNXiazT0QMgHcuZOw4f/NeU72/+g59HhwNfTh
clvJZdqb7ZqFlkg6vGBMZk+c89F+Z1ty1r2DqXLbAt95Tvn9ZhTn0Ktwsm4kQqYuZVSSXp318D3x
Wfh1s8ubi2uTNwmWUPWB+1VdHMeVJ02j6Vnf7Eo0k30DcXkSRWMFkj/tsV95E3dReST0Qa6sqfk2
TWCZZtVdKz4AguGk5NkPHVKMeGgK/xnwJxNU+q/kXEvKTekwFqEzROvSZP611VovegQJhqKiGq6j
nCmDjMS5e+pntw41xKHL40X+9MnsnBklgKYN6+vzk7ZISNyttkz4WgX8j0iFaGvPSl+LCPR74leD
/UHjlWWRCRMk4Zz6C3PxAMtdV+rP6LZ1AdaXXLaAZ2GlqfQ8RabetRaJsQ3G7bkqlisj6D5r/rcx
HABRp0+dxTTUCSpJ+V9Wk752kgohw06IBbXq0FdEDQwU9KsghmK4i3dYyk3U3nYJ2J5yNwhLppp0
dJaim76cB/TEQm9C82vzy20CZrpF0VAxQSN4aUd7RVYJVZktUXbQ/ZCPq4+cI3FilxHWu6lhjahy
am38fU6a5lDIt7hhuR+p+b4/i9epsP7bh+6oWPrpWDCDBdBDRAH2LhJyHGzckRk2LCVncJuQQ76h
4pkiRAXVTcAMPUksZLvBmFZAUbcDvLm0DUi2Bp07a5hqc8ty+9jIVp73P/2esF+n2jTBVbbv6JIw
vxi84OOznN26HIcswfWyEDeWdXZ61tUy2Kw878zmRu3rH02ykfB8CIdUPEoaymXyAFJx2vGCsnKB
yrmf0sbBYCr9cxMLlv7wzyWVzF74aOzqH/21J6kS35GtbCsCAxtDZiMWUCntFr7yPvcMP/ldG6/+
PydaQhxp6/MkIflLf3mWF88Qmf8vmNpXi0vWhrUJMfm1/FFgZw6tKttpM8jYdKxxPpLGrIUP6DrB
Zose5vXxreiM4AKm77AKy1rm9ksbJSLpW4O6AVoahip4KIQ29TTUJgxztmZBwkIJV5BjOp+i4dij
YyE7QcIlESz5p4l4sf+jZje1p+gzZQIP//K+lbrC2amfmLgJWJFXPjy3supy+3DSs4eqPol010k3
WT02LSr4JgHXqN8TrHFXV8IZxUb+LX/z2Z3kikGgWBvPKtP+qqIX5ChvVR09MKPr4JIYwcsSEezN
GapkayL4oUbBVvjNqsw0BHXK4A8RHrAuX2LtuWhWk2dQxVE3MNx+vo1bORU1xh/F2qvvpCI8cnEv
7iJDpYIG6uqott+lBd6WMCw7XcwEhkydqZapW2J7GNwOjbPy6rGWi5BrFhGpb88VAuRGWJGy3pOv
bmqWtQpPPDJxHGM0bD72fsAfYai6QC46xXqqpaIwutpuom1OHgbFnqMp+X/5+z8htwG/yuOp3MQa
yacba0cdOsuBimVtDcTKpTTbYWErd7t2efLDY8yP5oKaooMe/k3d0IytY7BJ2cTTy5Ft0Fw0w8E8
9QofRK6n1VYZBdPcbBnjXe6JSSdiqQ/wKappewc3MT9pbQyjmp6K0q92+cub+XOH3MJ5mB08VdVz
TSIW0hp46bsokJPIDjtiefIw4SN7jkC8e50evJuVD7YA5TcRwnlU8EzlSNWU+VoLy9+LUJBBy7V3
3OLo9aoappIRISq/GgJ8ykrg94ln3+xP/VzY8M1aCKLkoWfIZELTzfSFZPKu8H/PEIzP2gjdLBkC
lNRrL2ns2UtqHHLDE5C9hE/IiG8BDOV7Jqssk2ySEv0YF45z91W32G3ppWg/eSFt8amzFRhzYDFA
y+sng47SBTOweer4uuD+oASeraHjDTgkfRyBUH+WGi6f5sk5vABoJ9GESFeMhM/jdoDEjQNDUxbq
ggC+e3+K0U4YI+oenQ3o+8w66x3bjzLkgJiqgobPgzbWtxsr2WSYHqSHiNswo4g9xO6jLsHMmk8t
eUyv91YCVU0QQDoiTIeczEGLHjQ5PPnbXFulnv/EhbGfmSvTQI2mmcBSP2ngyJkwgOmv58qz4h3V
JxHS1+A9UgrdXLIP5dp+uCmYVa9Tqf8g0fGCc3Td+JhMn/wKtVLew5kDtTPB863XRa0eMGWzw7YU
CtL620yS24b0IgmRFs0r30xBg/mA3AlFhG3x3i23+6I9Vef8alm5jax2OJ1lVh5xFPNSbtvBSMF0
+mki5XBjF9Z/oXhsdb2dFJ27FdGLjlk8qQHETUdzL7EnbjC7fcol3vR88AE3DJn0Fi2l+rBaezsd
BDSdkzGYh4H0rmwic0X15twHdqyid/IQKqqNGzt7e079Cs6B0ZmXitSSjzxJKOOpP5F0iRk0SQLN
uQrE7fDo3DdBNNgz+ZE/4k2Fk4Y6/502tWbDBx3rFe5orezayh2qXuaNEBzyiSRPg4Ly+5dEhvoe
JItrkYilNURZCwM0aze73ukF5ndTJS2kCDFBs0I92x0JE4l4siHO3n7sM7Uy7mgSOjmJhquARJG1
VBGk5ttsFPy5vyj/rnH+rMEGcnQZFS2RRSq6m4qHLEwwcChGTiCSGBzjBezOHGFxLAiTc6g6KF7H
731Jb9Z+TT8zR36T6PHi/5hAFydmrQvhOPrNQO/jfWAjL2Y5Jgb9IGBJTvha1pKTWFy3rJZQxY91
khTHriU9CDjaTDoZ7OxUQDqQdiQ9M5fwWHhk4Zslu5Sr3PBimqiaOGE/K7fT5+t6+X3DCa7kkObZ
X6JDh8QgvJSeqvUzkHKbV5uNflyAdf0zOyJtFSdR2U0osVtmHXc/q0ytWft6dNWakn9B5U85pkFI
B9T427dCbJZdoSMnqYshS+tgsxaHl82LlpX+1NBFw6UUee7ZJ++rPhSNbHtsi09FJoHmALX6xvXD
ebu+dw681habGhHlD8CTvae0x/+DzVCqrsrx1CIV0mP3MOWWdJoRlw/OgU0jSLm1kbjSrdMHZOYh
a/Flj22HZdzywUymNbLf8AYWrenxbxdXH42BP1sY/GCdRXOF7gauYQzGA+GNWBvpQ458XnbM/eu0
7gQCCyT6UMKlG4uw8NewJG0UMLRfqkwTQ/k1SCDnFwEXzd3E07ByHXSVl/1NszMcXkGhEo6Bq8n0
8VlysmZcRNZEL7Lt9RrvFrBFV1mA07ul956lYJ3ZJRBlSy4zIfEQKUux/CEkPF/xMyFL8Bc6VES8
bbYtKdQcvBEGMgLCd9vjcDUGLxi4Rt4CC73S2dQCR0dWOymVT3baisqzmJvgBvF+fZys599Xv9pp
xQIDyWJDtngVxCCbeMamd/fEUi++XniZ22QQkLaXLPjy9FFngfEuzog1T6QASFg6unorK2CRwZsR
VNrs8fjcyTE/nVj/FdMfyFarVJbmTu329M8oq5mN/VnTe4RizSlDVsnIMnMeh/q96mML8fX+7IAY
PbmSnV1P5HIlMHOM52Q6EqcXGGeKGwsKbgpmPcCAl0h57Gt1aEWkfnVbsTKhyg+BJL/8cSGObB8Z
6wcHg5afwZNRiYZXX5B4M9lFI21ZkKkD0eRbzL2zl0M0yT7ts3JjaLBRp/VSPcDN0gphNrRWcXxf
fAKJxlAqc+3/Mnl7zSnZvsTSgONSRWPbFhtv5gY7YTkz29xUZ4JUm6ojN5JVi6Vp5dx8wN5hFRIl
b4PPt65ubwg3mHCvWdFxI2vHrxaxTshNPlj6OjLCHI5pcTnvM8FuZXzjpWKWanMCRUZFiBC3auEP
uYBajGUBCKZo2nhUGJzIRwhFwEUo4K3P/tM68Hi/LFMX82/a7hw1kTETVaZKo3ouPx4Rx5AZOax4
4eKywrLzAFPiYkizzCWmYa2OLybZTyqmhFBS0gdIfBXnmi2C+qlJsDsaYobB8WnZbpOckWPmD7WU
fJyIvLoWCRndFYD+yK7JG58Ebr2qGHzZBgl69ns5Id4L5XlCq8/A4J6jZfThjWMhLBWkE5qi2Rj+
hbg6WUCVt8l5FuUnJ5Y/xVNQZ7wNflNUljP0KmIK8Qa9VGBYYElvBx1szi0FXvzURc2FuDvakBau
WVQOAuGvgGYxX0GEd0mq3CHDAdhN2sH6vXmRnvdU0YqWCqHJe0NHEOvp4lq1H6J11cBVyhePyzzR
Zs/4uozmgv16lB8Mz0u4/gaE8cBZ09jFzX98ZTxcWtsYGApHoOiohFnFX1X3Di06PD3gdtgqVhey
PNer89SH7APbAykrgnhSElHkUJzM0cLs9zIvDLZz/6Wmxk4UU8h/md56NEcYUeveTIcdpiN/nOJY
iJK6GlhkMm1N3oEV7mYHVSY4F7xeGgxoTvIwLMXXsTSdP0WsuAioyPa2GCFHH53aEsmQB268wo5Y
+G7OKEoNrcGzARAec9Ozf0cbmqfqMTnJY46W0PyMFikWSBC5GlILbH4u5ZIJH3GNJ6HIxNWUyFNa
jFO+25ZaporNvMFQsEJmVsWGY92loMwFIhf+xKBzSBQcnCI1d8Yiu6yefT1U6HvuLOCqm+X8huLH
e00TNZASFaH8T9R5iWAcC6l9W60EtOrvoSJ2umu/Mg4+wfGrT9N694SphY/lh7VV4PF7w0zSEsyr
gEhcbzmeTXPlt4WPwVgPptZfpSjOA3O4okCIKrma2kUO4kFzT2WSePGwOMCGg4oEZBkZCUNpem9/
4E+TClD5+Ht/wn1iMWrv9UM3+lKM9IGTxg5k8brZFRHVkAslMoubh1OLDFQ3dqaNELqHwKdAWeaN
+2WBzJv5owrUiwOimQtJvNiVaVXhqOdXc2LvHC0D25oJtKNANYrjBXkX2Ul300W5jpj9U7bn1EzP
KkHhhnKXdNXT/LWleucy+SyK1x3cHKM0B7ydjp/6F1KszPq8qCYSzg7h+0H0nuyW2MDIB5nhNkeo
jP8vkPFzhttVshExzS1Q7J2OeVcoyyFSNOcaZ21CLmW7PKedwyGQQ+NxxlHMH30CwGRxLfbDEuYG
kamb1KMnsaSEl44xKUBUt4mopDgOUV6yfJJb+hqsoCMX5MBUS8V2a9I5vwT4yUo+9jbdBjLcyfwt
XYk0kH+FVOvhyfvmBtWU4eGTB8koKpk3HNmeGgTJsYMQIyvzTcFhrD0T9oZ1L7ScB7ieptK1uemr
K+S6JBp6c3X5f+ZnWabL5CxTp2yuwz43RpvtGg9dpU/cE1VPOJmwDU+/VJPbS+vSv6fqdvmzqnja
Dqj8/X7SXdckewM3Y/LYvGqNtyzm7/dC59kzfY5rcYL3IlCWPjXjz9ul5QYvKlGGilo0lUWZGPQV
r02HeRzIj/0htPw9EkEp+JTvRRJU7Srl63Se8ajVnOW+JwrK7Lee3WMT0APBrrUzkGxg5l3p8Kph
O49+UCesBbbINuiAPFHWH0KSGuymbFn1Jy6rXaakSvJx/gEptyvlOJcO3tdb/IHJPt25zMDkn62u
rjRvYAGNSS7oEbf2P32BNgb4jjJ7NinHgxWdelJWBVC/rKsVXkwd6OI+e19ZquiPwMJRkaAZ8wjj
Tq9rMx6uwzzOZmdO2hSXN7Z+ACRoelASLw1WdyoSWsDkKfjCJnTKbYf/L/jeYIiqU/L4t+eQ5YAQ
FRezHlZ3UdLsyWOCDf2ma6jtiejljd+mIJ791YocKTjtP6WxwT1k8BqlLON7wfPUO4hMcpfoUABu
enE+62O682fRLXRCYXFqtXEO8KkRJ6VyXCB8V5v9Lk1EaGTJX5PT1aU+z1ZIXWKThDsK2c8JrtCd
tlBeCHt/Hn4iBxirkahoGKiQ51GXHAQKbK8l0tfLs+jmArOWQ10EGWYjp2sOTwpmtIuh22yDBHeA
blV4zlqed2BRxkbxN6DlI1Zd7CHBiWo1yywSKPmqUa1tvarH5nw/5MZWbZAAzs4UeWla0uSHOnOp
5TevYexFTrSwdgEjH67zzWuXN+svgDDsiw/6nNBA0iZUYTjCX6ItFINrIBlEMSM6s7XmTvDsgwr6
M+Kn7R/hmstFY3uOcDPkm78CobqUPTCfOz2MVnTcDq9ydWkKPe1Cx9RhH7eW1P691ppRWyueOiS7
LjUBWBGz1sc0V3cZZ60Xjr/q0atOc2YKeApP1/UoXl7hJZhXc6yCQ62OfZZTLzLPRZaaFFRmDMRI
1poLrBaFDdtWwl/ga8v77FSNsGqFOiuqMxnuMt8Soe/bpjCmexv/mxgeTvY2xnpCPIcLWKxOwnFq
qEDrnZkwbO08wuoECWjJA94u6PKqql1CW+i7iYJEaWvfO6X4aawtnnscQdA4etN4YDAvZRnlswab
PmIvsOVUg9KNkynkpY6HeQszQ64MVigqsxhXivxnfefZshrBi72aklpTBiCwaL72B9XSbuQL7t5X
f+8OgUN5E3ES7ZHh0S55AQcAbZcPgyl/XIW5vh53AjdaHFM61R8MBjm0UJIqqlwDza6qDnAvFI7u
IPQk4mj4jxsmy3zbr1fH+p5kwKke5jQuAqhMW+r5aQBGv250erDlQFdvuH5QsahPqaw0490ZAJuT
dcJGs1DIQTQoEhRp1nXmZJ6arDeEMc3apBHU6KwaNBj/PmwpWXzmqoX+gx2WgPqBRn7wwnOq7aLo
Gh6IlwTf+0vNY6Z6PEYNESxqnYGpPl3cHfa5fjIu0SvH3ji32O/G7GWM/z53ShfWyVPmE8EtB3/m
h47SwxsMYasKbIInFnlRCcofusgtUAbpbyecOorpvo63XTWwyAPKKmgX8+32pbCMAsaNPXUrAwIJ
lSZGhurv2JivqMG9ZfegcSYdyftaKjA/k6weVJUEvUWPWLW+uUv/elLwfu/9cHN/ZQMzVDv3IVQM
idn7CjrxTKCPprRhbk18CX+vkOhO8qWTsjy0qm0FCGFFo8tpZBiiaa7wlLoTwFuiyRsGotgiRCvf
eUM811xWYwoMLj36Rrfl8ap+5h8/VkRzpY9+uIaNLVV/MbSG4autULT56OOOFx5XTBlmY4DnAIxC
hkFYoopU3zNEbFC9/4EZAeRSonaHZUd9Bjod7+SZ1yehcX5wG6bU9Pi8ieHlg58CpAblRfrP5iKR
RxWpoopCGrlw6Cx5SJYGdWTSPBaHcRCjxfbJQfSXhFulqrcfp3n2VaGrbHypx/Ywwv+7qyA2Yoz4
ftC6vL0I0TWG6J2lonQcLQEx7yIyHT2ld0yp42XxzY9uENQGvPzVAPykiyjUk76K26n2xA5LqPkI
IZ7CsEsZwzDdHZWoejAo/Kn3DJTorlFEb6OVDXKlsCSFhFdus+4xqN9mBCJSYG1TnmFNFN9YZsXp
sx2MkK6UJHcA64bwINJvmucfs8vr877mDdExqWpoKJH0nMsOLIz82+wP0rfB15wRkefSsVfrgqIm
FKErBhUyknQL9PmGx1JE/r8HiNptbreyu27H+DqmRH2LABTsaQfm7VU5QeelLQtFc1XDaIf/8nwd
CW9XTx0/iIHlIh0I6R5+SK4tfYnaYqIx5f4T7ZLDWxbecM2+IcRh7+UMkBjaWbN3VnwhmwnDsJmq
Ew4JYt7THpoFslK6KcJZUoXRj4EzmCvp+lYPUHw4ybmFeabCKAfD6NG1GfYknw9znEDIjfYraq8q
/IxCfelw8K0oXcMvw1gyOHDDS6EuyXY0iubwIMaOf4Vx+rKcqFGi4bQQrJlBFY2m3hb5ExnVnpG6
oii8JwdPYiFl6/McaaZMIW1/WVPaRwml+e0FAKpo/Ztacg+AD/zSyUHqo/KW8dDJNFfp4TCvCNN5
yqXAuoS/D1nKawLwQzfQBAN7FpkfuF6VXf7A/XJ3+8kA6g4clnEV+1DHKxBDZEjh+yFI1lQDt7C5
Co0b5LbST5MwhV4YS8c4mKXiJVRK1HI186jjdzxj9167pNGzlfseYN7AgUF36N9GrAHGCAHoZW5q
0BEomVQB8ssvpvskjT3Z5qu+LUOovWPeQAmisgZ7udvlt46RV3SAfcNuCj6VajRDwaIvk2K/bPBi
pM4nYM+01VGELRkkM1ARPrLO5zLXI6ZiauUnV8xF+dY05UBQrlfg9kk+J+Mi2zKum/L9OXsZ95g1
FwpUVNmjArF2D0jrt1QaC3ECPxOdUsoWDaXKk3wAWR+hsgxE6Jm4hvce/Um7jx0eaRWNHx1XrjHO
VsxSPJXL3bVDchgtSjQGGQqZj79Gkg4C0FMtucMHrN5wWQi2Y3QbnnMhvedvm/GWmMzVIcJ9EF26
7FP/V38D3PwzoG8ZvzJUYTobbZvDRHedKgojgbxHA+Q5z8Ba872NOjiLzr3hFhZiA7MYN7l6bjv7
SM2Tggwyyo0qNG9YobtSDixOm+pMGVnksLcBf/tLVvEFi2WCNvmpn3yDV9li/Yz9/LxyWMrIM5sQ
SwMtvW2bIkiWle8ORN9u669n7P9Kg0gEUcUDDbmo1/MR0urqwY3qwJqxxrwuvbaHqYCQxTMhERdl
RRmb7HGd1mpvvvn6m+NByEunB10xVHwZ7PS57DcQu3B1op6AL7b7l7bhvySooVr7vMn9TLMc7FTJ
3bjaca2zOtyTLru++I9LmvDaTcPp1JySSxCTmMEvPmBrLJv3q6I9agJ2ZwwdRbgnrRG7kMMzimrL
PqpPsVA4TiPVwafCzAj+iIEomuT9UJSmwnniR7S2nzb9bRujziyZ1m3Moio96+mqgXsaYxHNWYzn
ZJtyUH8U6rOcAV0m13HCw0TRmOdq5G247y/GFtl7Q3UQAObnfeOtG1x6hW1KK18DlSCHbNTfbwwi
XD5KYgwXXW5Y9jHQ9FiUxVZqbzTD/vjVNQKs0iv1dWuLw5rjRjwcGV+uCG+Wa9QipWuNUY3iN7BL
rOvVoulWpKWqJLSjVptlK9B5Hh2pZB6JCFQkd7omzVu5O/qabg6AZKKx6fpY9c6H8n6Az+jIo7I+
BFlpFf+FIeGDNn7Nt/OBQtA1mayWJLzyS26YaXhdWfN5yd+npQSEMVpHFLTpeje+nMGX7uVkbxqd
DjTM1OLFFzGxZuKiZds6VLuEWS51NIfusKADJhdPgy4ZQLdbQddamgWyaVBCdGdX8a0FK/JxnOTG
byGDkRREMD1eK6Z6AeOyQeoDzMqAC+6y58TKKVa4iUAbpS+JZc4HX4tdnW34ccHhQMMwdgTukgEM
e+AM1Afi3Hy8lWGdJ/FJehN3EW1MdfZoS0juO7Td7YwXQC2eX66JooUgYPMxUbMo4bLkEX+Fxbyq
maWeb0v9np+QXGvEJjpqrXuNEBZtKcVaPhtvZD4BQEHgBbJdASAzST9dDR2Ie2TayMpTOcpAbenn
cXmzWXjmgWfO9U8yM/L8xUAKhDrR5tZmQ/2lW4LJTPKIvabK+KHe+vOkT/MTUyEN7mVn5ZE0uKgi
H/afqdJPBQZr5aS6+njzL4O1jH/YXRHJxGFqPM2tjUVzSmXBtPgmNGtMOAP8avX51ZYWBKWJbrWZ
quZtr/sCWDkEalsUuNd/e8r/j7YQKL57IIdqF0eLu0VqtMkEdk3dZhRcaj2fAA0jRK89Uiw4HODi
25JYXe6ZqSSvVA4Y55472Iyh+MSSgFm2faPGuPUZpWYtY+6OhmQ1b42o6qpJLjLn+T6Di0hNf2FK
0ufHL2CTjBIWsOl8zafhykfwkw7xhfs9DOOMjHD9/6Ed+AfZV63BLm/QUtOL0siGri+nuGmujPbx
uHE6B7Bdk4+q5plvj9gIrePHzCn3FRj+fxTNidnZOOzfZ3c8hxN4WoBoggchF6/rySjd8360x6ly
TmkrZb/uhrho0Rq69qO+RQ1sh/YLGvJtImXJAauYri4yFUiomRWQ+mNB2dxUOoPHANwpG2PvQfEl
kWaCNiDtCYJK0JfzYyKTs65jY6CRW4RmO0latVHSPI7oW2GWKeuQ2iWJwqokk14mkVXISULcuMLq
5BsqJHH6ots7Z+P8G58aWMEqnv2tzrXvBSyoJGAYw4B0GGIDgF0qXeMe6tXWjZZ9dmNP5FFypa+p
5sHKxLicG63WrA3bQQ8NpuCLBp+gIVhBxnCWGoUiDPDZCBnE4WRjPMi/jVOgU7OS4w4lP841HBtS
T10T5mGWnFDPSDm+jDqD9bouW2QA3ZQ93/EfTIKJN3/YhTSRhUxa6L1c24fWb5IjarBel9l0r1a1
1ChGddslpsVtmhTiCQoMnnSJATxV1wxF/EBmmxd86I3WH2vlTLeIBKFylV+R6LMfG7tcEZQZfUtU
kPd9Mdu/DfcZJP97fjIInrxgZFvO0TF2zreJio7xNeZiKbvfAIgLlUFOT5pneRo4bzmcUFbF4bhp
zVudp5/3xUMoFZBlNFLu7ZcVWXwUkY6TggenJHx1w/R8luzPTC4r5d05RLfqnEZzf3nLfOq0bhJ1
nwp0K39aJn02iP2p/oG2h7CspsKyKARm65b5GWGS8fRW2Xiia8mio2wr37Fs+hKp2shIdt225PJA
dNKySQ0DbsaTMZSbXl0nI33m0hSAlxOkSbhof9k1pZ5KUTQP1OchyvzkRJa+ICeAY2c/Ctx5n0ro
UYK4+x9qrvdhuy28Q1WREpvH4LCkuH+WM/LJerH4KrO6jgrgyNRyyje2+y6OCqoPr7+RGQZqA5eq
yLlx/sAtPvnrR+afTp2mjCduzsn313CmXZ/00k64LqahHybhtV1udBXvbKJNv8poqncvinFZH/ih
nRYhniGsU62/tus+qetkiJZKIHg7xYRPBgn6YDYYHOxKTEZEUU6+KuL4MW3oQzYNu7uGR3aaJOyM
8zXdVWJ5JJ8jrrw8YRBVvLdtP3MqAcpWcasXTg28mwPJKmVC0xrYwOdMuwFXBKqsUCIs+KNMyCtG
kaesjtMeIOL4NoSTeT2PvMFuqE9lNJcTqr1WlsfoObGSTMr2iyUjd/zoR5RYW0XJHAimZ6IJ25ME
GXzXwP+95kKH6C7G8cegJ3RQ0aiEGZzlJK6UyWQVgFPQLSp2DION7HaNP06hB3prB++AKzZuoGDA
4vpJJRLTKzTeXslMsi1pz4Zo1GlpQiSDuKgaBFJ6xxKrwJBcH0Q0wHzqlAG1Wyl1FXMtKeO5ZrEF
L1mBlcRTnY/OLHaHSsMQwTdjLnQQItKvs55P1LYsoSrPrshLIp1A8gkvLK3YcC5v0luQN5RgIqAY
IeQ+xjiw3Jg8rHxO7OeDFNX9+FZaFqSs18CfnidGnO3UXBVgJDFFkqTD2/+qa0pTsKk3Fo/uQV55
vmSrBKjmeT2o6su6YTCBHF+F3ctlc+GA/PQ69F/CZoABtd62re6LyoQfJtUL1yWch7yDWgbCwsWS
IC15S9lmicm+jfDCShSmBkGuY+EfhTFjJjy6p6QYcKDLqZqhr0ZN/6vnQM3aGXvxKOCWjYvbQwt2
sU0hQ4O8BL9/8+klAqvlhpuMfftGCVjtzsm48tYLxG9bbDIWt5AsionVT2acMeRT1gdOwmSqKVJ4
QHQMVVs7spgFg101EHxpesnojleONcmgGhgiBGuhtevylC2N3bha8UNC3Tc7FMd0vduwcwvDnjU1
VLws9iCOrWJUV2mKt4ALz23u+QRSaPjw1PfXpc67CAblPBjTJHjEsMCfIFGEd72bGc5s1LOo3/HU
BL0aANLy3Uab7ijsJJV/Db2MuEWw4tgQw9JmXq7Ro2AQG7/iZ6uMyaVMZiDpP1FWcm4wUYyHpeTn
PdwJSjuGXO/rXznoZrQnRrrULavmwS+GBF51FSG8FhZTQ4mIbBh/aZ+d9eCKGF8E1NtW6HpfV3UC
xV2n2jCe13opJ7KryI0BFv6YxLA8t49Yq4fXsElRroWaddfUIXsj1d3ECf9Zmm+B+LTqreNKomos
z49EokGigmE7E8oUiGWDKDqrYvus+X4gqEYRUPuyWsMSSTr111DHiBfY6MocHqAytIQV473Br7E1
QiY16R+ekwh0WB+3DkGMupmX7vPwqpDu7dj46KSl8bk2uyC5elGDjhiFX6lWchO4PuiM1an5Jbc0
kb7/247u/Xq2QSZ2HuMz8p4/qAuyxtIlrOvs1B1jg7G0H88QtsRigUZS3T0CJ23qtwNBe6ad8yK0
hGTM9ZlupFpMKhWtzptEmfrL8rfJ9Kzz+8DT1d/BLAKIFlE0IiJLV2N8f3yTLFGoLln1B66C4zle
V01pcmrbomPZ54OznmnQUJdNpV10+w0Tvi5JO9aMqt7x7acduFXmBMwH9p3dylpRaI9EaSTeetoj
GA6Zro9QWg8YjJW3vfB3lF4RipiIl5InQNcfy0LMz4Jnqhw6u14uqedgQxVKOaj37O6CLvFAgFTd
wUHSVx9bE3/eLfDvXxLYVkiKqurMt3RjKFu2vDCrAFn6A1OUrab9mM94Enjny+R2gWO7imQlSvQf
01GJbnjr/Vp6lGegJFdp4H+u8aRQTRG1yqq4fBhym2WOhwAhPXI4arZmKZAsuPUZy+/jbvH59hF1
vhfwV4S/+IHuRlcrggsC5WA6GUQnUumdZA9J6DiYPaUuzYoFFBDghqhBij6lO2mbphrTARzpOAqP
jUkp8kPZZY6JVpE2AAZlxpsJ94nKk/tOWPEZtrZo6IHz1f70nbrbwB5ZvVpVmvORKGyWvY5XQhGM
jxSc+bta73TNW0trJ8Une+EOHvN1yB2bT2lE+H7kaFzRp78FRZmXOix0h9AqmzHWWfQ0PsBRG1sa
bC7ixE8FJKbGehnMRge6rao6KSS7gxbQ4E6oWVjVLE3LYTs6hsth1YySkUmsDvYmWRGETafX3JEj
iBcoUJLmtBdsJRt7e87sMCgi83Nrwuj5PVFDZ9jD9+4C1u+VsoI1ArRlGAvJUFvEM0+hNQdrdxJn
BBVEgbZjdApoitQfWyb2Vnae4CRLB8d85yDSDzHnR7J6EeR06SRvvsBnHWpm2o568AA0N4NTiXhd
rdvn+Ek6Xm5Cu8CT/K8EIAr5cazgc6S+cpTOef6KR85lLxQ2PVhiITFYF7IFP/8rCwkas5sFj0kh
WHexnWHyc7W1Z9IWfxy4r9bXjHXzumJXvU5g4dGTO04dGlcbKop0U2dulNOKhJe+q6RDaL9GwuhU
h2auN2wDK4VsNLWU316HX1SatiuC+C2gIn2aPGcKhspyujaO2ddfRXtf9PWgxWg0tzgB+lPMczqS
2G/LGjcKvL+0YUF/cUxwzhKZs2mmLFQhtWbDoLIaVTU2NSU4+hpsuu+QGRfT8iAZtTUH6Y0wdOBB
vTVWYJHWbS9QytP3Mrb3+B922G8TWnKEGdFjZvNbeRsiPTiWeFfIluyGF8nwfjuWkq+GyOwpIcP2
2g/ZDP0hDgDxRffl5MO/iU4ysEMxvdcAtWOCYk5E0NYdmVBOXDia2h6QsOsAuJ9Jl8bAlgs9uKzQ
OzJT5rciD6DdoN++EGU0BM/VdqPYCfiGSFVhz8sLSfAualJAz8kJZsgF+Ho1H8f+gd+0py6HXfuM
IyN/C5LRLRxJd3Igy6tVZ99S9ApnL6MPtZhFgrrh0nnmlyBQp0K1gIEQ1b1Df1fs9gBrW0psjc+l
RrJNjx0HJQHTo33sK+J/3Io18r9Z4ivF3bsADd5tv17Pm9YOVAN1poQqHGtfy1xDuJ0ZXlUQK/XX
5Sqy0dpvCQq0ST4RQ6mnkbeC9xMAjS0IDc8huad05Q1zFABTuTKOlRLMiTle8LYFIdRg8C6vSDru
aBYCpt3FqTu0jJv+Q/SjmLOxl1Unc7pgtKlHNU2ZIqMRdGAkcpqRwxsFPkRmdE19ekd14PsU/jll
5XViWiUtD8XR1lNPD7fISA5uKBpdQffDu1j5L/KogsTSQdCfxYj3e0DbURE9PScbbeRgdaRDbpQM
T3GVJ0nhjdk0rY/AwyScVP84voHLs3St597zXWv1M2OlHDnUh48KaRX1BwNLhgM6RifP07SiK3bf
i0nOdQg3gDzf2ZBOHa21R8fRzOkjlh12c+FzvAu0G04n5Px6Ag/VzXAuwi2LPWizb2Cykti+MXC2
SIVbLDQnK3FTMaMb1Gbce3yjwMp31DDq0/R8LsqTlURQaOJwJp8myJ/I4/Cnryq/zKAAGcUnmil7
pg4rUYw4Ok+QUqgS5/INK1grI+FQ1vvP0kpwlZSIjNRIZIugBFpe5KyLWnJHaDLCgrWuHw04rKW5
hMzxG4T4vxu6qVN8bpzvFZbwa7ijP9nKbz/FuFjlWXb5QI5bSnzvclU+VS6t+KfOGDURgbwYqAs/
S2coPGyFQqj4YsEEMgj/g7DSfNrkd92sTlQ4q1SriWpaiK4kQ9Z1Vj/BhfAHAJGSzoDcOxnBwRGB
Z82jTbXEMNanf0VNWU8X154at3GLVyW7ZABpwXJWWRKtZ6Yy/bFec8nCe3Tgr4JkUPTqwKvcK7cr
y5NGbwSpKzxXeyENJSGE+pcZe3yI9Cyoys8R45dmvM9YrE6eLO2MwNGpjjL1TvZMg11pETwCCP5r
1duJ3cFNZLAVc8TXCdJZ+oe+29NJo6WPHJfQWRoVbNDB0SwA2OcAcU8IddF3hDW8G0d2iu1e1Mnn
FSmj9ZohfREJnedSYw9DHTl+U/p3cjF48eJCdkOKz45ilORXUkBSwlhA5u8wRKNzvvgb0Fvwfbl/
hZyYoa3PVaSzDyi9+ani34uFi3kuaTIpEgBXqbVoIH2ZKt5Q+QdspruMc2GmlserdVJtkMG2ITJU
P0IspSsqJFUyjUs6Mto5JPngf7KOt2L5M9oFGA+IYzwt2qnGW5r4hukmdHTR3/UYBcqI0UyYAl5E
ikZXv3x++kKDLxLt0yaqf0DIwLFg5Dpo4RIoQl3mfJXawDo3MlV3Tq1KxgalmsF86kFXTANb48Zy
9NEwV6MmJPzA2CPiYJzrSBYnozZVRVOHwx6HqnRhiba4cm8FeaTwDEOLxld3Al0ZRh5FH5u0LR9O
ckDmDzPQCxW2ZmliW/h1DxwlxZHy04HRoqbqkqS4yfKk3cnmojRcvlTbyrgDZ8tzABrLlvcyBRch
KE9FnahxWD6bz8Tf8FkY7ugF3/WMVVc+TlBLXePxTHowGxu+QtlngHSicM1RVrldzQUGAy4UqLfu
RHbqQNSwLYMO5WlfcoQYyp7DZOL9JohB5TZyaG2Hlxd6whAn7jdJnSNcBAIjCWAAZhJYNf39UPnf
16QwPpAcW/MlmH9oTGOukm1aKGm4ohcOm1SnoeMaFyrCltJjQ5rbzSK8XRAxoQukLVJ6kcoAJHmr
rOpr4Py/xDmBsfnfK60TgX/WN8b5L4Eg8TvV5No51ssvw3BnqFSesSVV5fZQT0wUV7u8hvfnRBvT
SpRo+ye7ttl/+flMFYodQ8bovOgblyntgQQ65Bkgpgm1qARxdFMvDaxc8i60GYLrJUv0ahA3z4MP
OImT8lkhEO8kVjSEkqM0w2Gi6Rh5w5fNkMZPO40CViyFA7SLeQN9ppMfCzej88ADmtlgCryxyFnC
c3wwAwBqBBTUi0oGTbrJq5EsXdM2hFyE7UvcinVc7YhGUMZbiEwSTZ4WaBN+kFaLe0RzS4KS45fz
vMtaAhqpwTftuVaAM59/tz/UDRWCFo8y/VxDEso/i74WhLcbrDaFlvH2nEoe45juDhsgWGnyJb0X
nqvgwm9SBlzaMbMr4Tf82hdnisBdxyV4oIXuDNjSxDwVsuhiv4VQcAUjxcMca+jcQOqk6LKEkQcs
QGyOPpAEQSYnWhuCWAmFoU+NxokYy3XtzCnW4OW+BU26pu+ZRk5rCXB3vkfT1NFAi4lTd9ggQsQL
a/QNyM0DJ7du2zTVnoJSqOmuS6feY2bNbMoz+aBYhaIVEAVWlIpRV+Q2Lal6KPTdGOM1btVoo2Bg
IvJJ7rJKMXGGSim3as64CqvU+Qbog0De8untSyYU5/0By8/2lctesVVny2lgQ4F/9alJJteV2Uhs
7Sq/fq7N4TsQtknB7udFgN379LJ8IxNnxkZCtKTQRcd2z3q8LUriQTcgReRfVO7OfI2tPCMxpN0v
MfYxJDcrdL/++tAIWueH2xWqYP/i8uQFre5KwEk5W5eZhS9drvLqlyXGYsJ3ISHmNxccjqzr1Pyy
nM46yfTPrP5stJefan95NUXyEHL/6tuTuNAWmNbEfKQ9SKf6/TmjQJjkNdHqylg80T5ABeLwKwYS
7WZfQKJiQOhcLKUw8yLmIz7Y1sj7RZT5iOwc1DvbJ4t5fqOdai0KmS0oq9I4JnqyOZ+BqF35XfS6
d3ZEHJ4mMVWtnqdbj+EQfBVsBsb/Y027lRV21Bg8HGxou0uZPxOzf7QhvYx7L+LA48GawBPv0QWK
ILI7m4giWdsikYOyJcD691cQYPzM2AGD/UUoicVMjmVc9FYDbZRgLkzqzArT0VfGQYa8vIeAPnY4
lkKmU4KYLeXJXyCfomiP/SJjElfE4YnvAA4FbX3q+9pDL+kYEyPCnMU81b9Lod5n69gxrIP3B7bH
xxcmGYCECs9nYSRDkoPnmfsq06anjR4IMG82kH9TtH3IPdyMuyH+igSXRAK5chWjLhOie2nif6Qt
yVHUdl6LrTup0CjcH8af5dK3q3NCe6adZ8hCbo0RV0j8Qc7p0UIAoYL72P8Ipq/fbo/za/IU7Emt
CPxTaDR0WAu1bbmGU+XXmTiuemRXd6fHQWyXb49OS5CXXmi2gW8ikhDwpGHeY+iVXS8B0HbAMDih
+s2dRMO07sJMFSFNamJp2X886zwaUuWFSlfWuyU1Thb8ZSvEmpjHSuzL1HfUgIo8H9xe4SpCo0qz
ODFvbLLsdpCYP1kHGuRlyp7UPCXBuQqTqcRoD3ZhOM9nWw7Hy/RehBQC13RnP23cGPDCyzGuqV0v
tqBT48Nd4PnLg3BoQTWkMISsaVAoqlGcCtlGZxshbXQZqGsJxwfoy99GZzJuTQcvAmxzeLKKIdry
eYYQ5PNnUp+4oP+jo2mzHxPMGU0Ivg6aA3nO1E4uG+Qqxv2ljwRYRYPc1mzAbdFyyQ2n5vKTFeuI
/SGVfA7mOE0P43YeElpK7Z2IFtJFE/Pz6TQf8vQHGKk1+u0GrRdW3SpiBgP5fEqvwwJbbHfWkA/p
iwZvdIxB7IixRT8v5kWml2Yk1Riii9bQ1ZDN3vHLYu9nKz2ccATJ3UdHgEgDaeyu/I0TrMNr2PPz
GGA7bYC8lHy0nwMp15nkzh71nRvwdLU8uNGumWy1PBiXwHcsUzjd9XcFXhN1mNpoXttJ0goWLRSZ
FCGKIwhQe7t7D+1IswBljnq3qKxq37t72QOPPnYLD31U0nqpab5iaD7jOfRFmiIq3nj3hWKTg3ND
oAsQ+1y4vZJ8WVXcSACrzgzq4/ODBUC9A9/9O2oO2gpULOXFTxBtdDhyiQqIpDkIU6VAXmvwUfxg
FWzCf2MsnqPbBGNULwb4AB7xq3AJMeQUQVv2wL4WPw5+bca0sQOK6aMjlYxK238lWsT6eV1czyd3
u+LrEGkm2EJumRuaznt+XO986KE40udNWD5oX2uJmMjuEGhkgUfIxuv44O4KfCuTMjBxxi+hxmpJ
OfvBk1Sgd3p+SfjbOTXAY5DrTmChmEzw00hY4qa+mIaqtJlOVr+8txkQUAQPiYhuNd+cZpCXU0Su
Ld0fDMNt/Vo7ht4gCDJdqyH1c8FMjit+0ifTIlVFhrbtkmYhJR8inJJpHEVoezXizI5u/4v3YHZ9
IAzKdGHAvLjucwzLUqq5Th3j0lU2tSjxPnYXJoDYhWsS8/QwkfGBuwhT1VbEF8x98yMHZGl0cGOg
mQGE913GLUFO1e61rhhPOY/P9Ps3Wpe8bDRd5/fuuoXme1tm8cfZUnGYduWQJNAJXzIEZ7DFzwqM
Nt5ZHQY9TyI/ULLl76Fb/NThxkRskEkss9hbfoFerUxp4d0wKM6lKjiEWjhUEMRIIWm2ONgNEjFv
8/fVxPEoolBKqsATAqiPIjFCjOQ6vwXuOJlTmjGn7U0kzgAjivJgSqGTUvzqbL3V40EDPpWi1299
mswedcI+GzQJJMIxYWOORKRJeetd8tutvfChQ5bYO3WAfyhhxnhZD06M5rHhVuk0zqaF8B04X6dP
AOBILQRQnJ9ps5qT8eAZsaUKcrvWcj2ALjBFMQvDzvU/FcJGihGo8MsDRV1XWRscPTKAmNlUXTO2
G2DihudakY8mUzkjoBsscUP3hrXngP80DaXwG7/9Z3n4HehW0E4orT9kOJ1RcYCzJ7kqT2Mu16Qi
WH+WLcpxeNBSzjEuittFyJMf0z7jDfHHJzZqokCx40WE98afLxUWl7rUsDFfEohfpaf5Yh1fMkZh
ofmlLCtmsQTNTbr5RP77KbFx9lmuzrBNHxTWO9I7D5CUNEbPtBlSv0thwhxeBih8ZGLOjCh/D8DD
n1pxmYjuE4nz6hpFrPAQxJP3Kuy9h2fdllO1reG2ulTZ1R37iGGlqWsNomHHDRRK2YcJigK25v9v
bFw/lOOvzHZKwK9oN7Cu9tWz25EzYxYRB9Fw+eNqiCIe5r2yRtMZMapS+L8Y/W3lR1MDLPXlluAp
d59J7JS62nrNYnDYSkOyJvMJlVtsKzr1RyzxsSL7x46iso34DrUgorGmNNO7p2DE7VuiBH7CU+oc
8qOn/FmpuvTfBCVl/Y3USC1MfckTfpv7cfmAoaHh6tYi7FP3Kn2+HbpFSi1ncMEy5vQP4mkxAn+f
WmZ00B0t2TZa/KG4Zs6ZrjESbazLvOUpEGsjIarnA83NpnrHEdyQP62zz0CV9NO11rryL8PasoHv
TZI8mQQt9Lvl17tfjAUuhxOAfUORzCB4SflhZcyg7xwS3uYEsrBkdwnGH8yA2krHKc//QQd1RwgD
fj1eQdA+Lsj0rudgPQh+JQeMwUG4K8zPDxeCbrVLs0P8nqwNE50M+hnxjM8H1Mpu14tVL1kxI7XA
2npLeubNV+vyVxhAtZQuEi3lp6Nt7O3KckWMzGzLtOI7ynFqgYOKn43bmx+1e8UVp+yO73JvRO0j
sSvq3c01ViZ68znrb7WOeQ1cR2IakLwlrK96rPWSilHJg9NTCmU5pCp9IovSUuFYKszCqsMNsM/p
5gLEc3sKGHhXeY9criWaruS3/JDur5ALYWU35GGJa+KIRdem+xeiqydSeI0se8ewuWDvG27OedRW
M5fWuobpinExxd/zY7TX70UfC1S/OXve7ufOJ2q1ZHfZAtdjxSkbdkMoUc4cs3RNhRtcM+L01W2q
Ow5NRbuzDe9c6F0G9PFdJZV5AWvOfhpOTiil117vhk8EGiShcvUfRJPiNN2YLcn6/NdENfCsImXv
zfiA6jJsgKW7UXL1aDgwsyA3eLXl7rwDIeGmrJJs46sw6p67nH+Vtm4I2gMmCOdB0rLDel0sw2zK
P9QbDxWmXgjpVZWmZI1Mg6LutrLe/lL/m9+Ji7l64+a2tLTpxDDR5U4RO3ShZY/P9ZeEnadbHCkv
WArHDdnK59XaYRLM3L1s5B9AEPaN3LpIKk3lPbzhueKn9Cp2FLbsjtaEGT2MUKStr5lF8o15dpSV
eWLq99boDoIDqXOW2he9FTNauQ8tsed/XotZB5OHtqvRUAtLDFro0gAFavNYSrwpHQnSwv4NmWFb
JHCdVxFF/xK5cRmm8iv14JWKcNfbOBtANV/w4MHErqmlgs3tEaF5IQ+zVOAfX9JtqD85dWmHyp1F
vmmPfYsxCPbhlexxWwB61VtAAXe5YPX5bXgmmobZetnehOrzwObZKhJSWnBWDyf0jZIZv1lLj2ac
UFc6VOOX6qNpfSnZUBZOWgOuqIQ09Qwjvm/MBZesE+iIGIsWPpZZ6H+enQC3Gm7To4qVzduCY8YP
M0exr9J35qJ/qMd4vB97CSBsXeJPqWy4AMv5n43rg9y4sMk5s2uwwr0RfF1Ys/G03muuHAcIpO9r
IUMfJ4la0FONrKwkML6K/+brwONDb4Vj8xEz+siXqZX5ILYuxhwqkGfCsKHIQ6jtW5Cm+14LXR/s
Jc2h22ibd6QVbSUjDTbwTwQ21RV0dlvB6WLcUh/jXb6Uhc4ZFgcbfKAxYBNMQUxsyWjyQ6stOxZ9
UYoIbZPtAu+2CPz02QpiJq8ugRPpiqJ9Rs84UlZIs+eZvLtNYjH32w8U8g7kborFIrdVV4wN4cDR
VUpt/HHpHdrxKy3MsQ8UTdriH4NIQmmlh5Xmny9r1NS6pnQ2HlG4t9qVNRgHb/xrVxmBr9pi+Klw
PO/7ZaJRc0wYEXIA41GFshSe49j3Cp2gZQuRPbxZj6cij+BBaHvnyX76a1meFHTFIrhOf3c7Q39h
zmkRMbRJdkWEJOb2p4+TWo0Rb4FDJvW8zEJVl4W87XJFGvSkbJkmANk8wOYXmgNCjqjRwVGXYblA
rsZifMlpgHhZaCkco2f90u5KB7immUHG287tWYLjhdp/NwBKYXkG48ir2x2SI+x4Je8g3FQm6wEQ
cVgIYthQj2WqtDb3v3esbRFQXVKh9J7BsPaLAeN4A515nbuwK8CRF59DsfvvGBUUo1SzXt4Q0tuB
wbtrvbZjAungRmlSOGMl0bVG8YLdddZPrKmVvxUrBzHymN2H/qJFu0u9qjy4f/rKwI1g40We8Y1x
daf2dFmB3UNutK3aDwELy4XEwhI3M3lhEM7LNBFT9Yl3PjkrMzbx/xz4u2d+7vXYwbg150vsSdSw
zKameANjokYKH50GXfe8g8SttphwM3JKFUTFpPipoIRlWv5rwcCtKm9ftDopwPGVvIx4Xy8LwFPP
BSkYcCCFvLJIIzjcEbkGvuMk6l2iePnx06hNQwQohTSCxzPYtEGJsAz1rlKe0CQ6fHkoNL1aqveK
/Q9dgAyfCdoO1VckIXTvQdT/uEBIaaq8kNK8DcZ5Cv/LLDqg/CWd/3vW41V7IqmokJXXWnhEbtsI
wshjWPaoKC5JX5rZT7ObWTENoKhVBvbt7B3CGCpk5pmHA1ZiTeH7nPNRau1g2jhV1Ym4E/ZnUpED
HdbJif896YxEYdETIuZGMMWb07xEtnR0jnmNbwc3yFH9yjNR6BTsUrFTCjCk6ItrBKX2C9QaElJK
jzm2j9/pKhUM2SmF1W0J5G5JGz9RVcj1okW6rTmwRz6HIhe/Y/wmcI5v6hppu5FjJ5q+ZGQIrXlM
RuPP132cSeFmMDaytU+zgVVTHBerBHdpadHPLQmZrZ669iDj000r2ARQL+pg3AA17K3sL8DyeY/L
dlXphM6+FJeYfKLS5BzF3kIs85+nOSA6hQg8ngj/eccKsH+Bu5xHZCAc3KvQEXaRGAGZQoF8wa8l
fKpnVhgIXTW9eRyGQw32NSYoV+236DdjzQy0KMR9odZ5IhFjLAQNU25oNu/h4pz9udGJsemxrcAO
j5uXWPq14PvBirvgiQSIaIetAo9bk7XtsHXRJSgww1m81zm93Qv+3uBaPkLHRz0agC66IO12Y3UJ
0Lm52m7Hy8gdWDbRNups9kEiJXbzZfdsFUldwUDOjnLvhvD4oRNg/H4pjm1RtsEqExZIpWuKHnX/
wQSTzzPtcsZBSNWH7+LMlucohrQlo/VR4yPRnk6ga+4pQB4RIFoOAuXdd3quMt38MTmJ9i7jVKvm
ZvoT5IBE6ATYEQLpgkc1XP9G/5oeFS3Yw2iYNGDg2SShBFucpsynkHndkIcntnpmL8GjJtwfbpxB
M4gHfECIBr2aFhRWXpO6ZY/UZbO/q/6QvWHcXWjqBms4rkPGAs2KO/UabplJaOJMB2PiJrXggT7G
CdSU8/AX5BkDlMAaRt3xeZRGNE8y+mxPiIynVym9zsRAxgqzQfK9voDQBlhMRsmQWXv7d0mnhJ5N
gWr2ocMRdYu4t6wjwrH+KV3CK66TcroK5Owi15jDtN9MpCwJ7QI9ra4y8uOOFd2KVkzRVlDKbVTR
PJmWRqyvdTZKdywPXqOxMWLv20swgWgIvDaPcFbSP/qTsLqY+qS1PHpMHrwM6+utWNCdPeK7vjZ4
M/NnJyUcUBeaBDU+Dvy20sekXdIYV2NVoBCU0Enkxc4fe34hVD6mX+zJcQ79mHs/PLfSp2v4t1Zs
fuLWdT47C60WvoXWSp3AblxGtc3q/ErL0QMxaV4xyO6ZJFvKhPSYdoSvdEES6ahMxm5Sh/czftDR
uOUruT0ZBXNSCcPGKSALd6aPDOVWjgIQs8aLnK+7ivYHPt1dcw9oeL0seRveKrOne816jR6Puk4o
A/sityOcXYZAvhTlGgOYYlEXgKEEjv3CWQqMdDuXfKU+4tfvm/WTanTy5sEMtgFuAXhyQ0Nnbz4b
SUsDjEJAgjisO/urbpda3yIuWu7pKT0hSztmzMe18anDUOU9QiQW/odJoynEvkvm8FygVurLdCSF
nxB0nvqw5VKiEIRlSbyuQ164M3ZxrIJItagK45eqgklE6gdzgqrZSyebI7f4jzyhC/eohMfp78+F
lrmo5CXEnUnmd71GS2wycO7W/O4qO972ZNUWBJowpqiVuqHEESujrWZ8dUviwLH+CIrn2zQTjpaj
yT8s/hg63HKiKfTJK2Qyn2TZS4Dwz8xIZZKFCFEEUFmBY2j3paaIfxQggnhcOxfR6Xmg4BE4fDT3
NMlpLzeTfz6PwE6Bb4/MD9tNim1JkaZ6H50OOZrulbxdF3zWTz8hLM75wDTw6j4HMnbJQO7GPd2h
jfDTDWTb3WSonAj9RnOMJGzyolB+JCtlz/1Tjy+vYO8NIwElpzn6qmfWySAz1RxtgE/eZPFPyHNI
kamVRjhgWGtii/9CU4QQiElHHbCcfeGYdrTJemvPTHocZvuIEds4TaMX9wyxGLt8Fol51UqJGgDp
irjLZK0fPJm4CBluoB5ZJi7l4HxOo/WMJSPMMKmEHApiQR/a6tgQHx5Fb5BM+pkIgTiwyYnPY/KE
jD8LPGRTAMuScbliYSYw3PH96KQ1tvqTtdmpDnGqaRl0Kfgz8QWd+yscNV7GAPUvwKC58fWuwiUn
oGxSVHQ/3J+8eytcoATHP2dDQZJGfD/sb8CAP9fC3mXkIooOB7RryAlEnz7I+Ziawck05hBWm+dj
X43yfcSJSwkkkMS7hnPQZEHbkwPxF4XAlJYSGpAkTCX01koO7beHw0WmN4G5Ixkqn7qA18CfKQ4s
6qkEjr8aV4aodcFm2YG2o527ige58lTanqX0n+odFpYZXL7SAEXt6KLx4W74zEVsjQCD7snyFds8
o3i3Ypz3tKemI3v5tCsSBcWt2dza8W6fVjZL0z2LiTRsH9j4izuKEmZhhtwpccc6tbxMujMRB0zJ
roNIHuFWV4lDIfXEmlXKCtl0RaRIRrN1NbLbVoyVeoVCX/tGkjqX6LligUgBigjl59q6K7S1cgwQ
pXlX0sCOnRx/cnNWQ2YlidzdQ3T566PwtAY7x/dW3OOaNWzauWSAp7URb6atlVsoPWxJfIqZG2D6
3tTQu9bBr/D4q5s0hi2/P2I8PG7O7sBVyXQpo0tSGHtJmPGRl18lbOt9MXj7pTBI9nOaL+WfOmn+
x5mgctW0ws7Fsk+v27WCxXfz/JwC/1eSESF931thhAZ6e5iqvdpwrPmVPPWYpApRnp5DtMH0T3dY
K2yQ5EgXbH8JGXa3398/MTi9i1K+I78cT3+mpJ1q5HNDbAZjqnLj9jSUIfEZr8WKMm6EzKA4fhJ0
kSNhMV+uetXKJ78Jou3knaXQWoTxSLt1wiTqTOx6zgDwob8U5DlbopzCU67NsYY28XMuvXLnxt9V
e3W9OMr1RosUWDKG4OXMfRFuUh1b0RSFcC6WbdlyVEUZnAG6rwxxarhT+nInkv+GmfX0hAKS47Io
9Qs3ZIGMTUpP+6YBVJ+oipRCf02W8cJ7rnkyEA6YmwPR6QlnRT2wm55ChUPfUDZAzYueCd04gYje
Vng2lBkTEZNzNCS260QmI4Yw1j7IcG4h8Kgd0CePcvaHbaPg7RSIrYacrnfrwMw8sj7FG+DV6ABd
VLBximiFoaf3i4l+jBtphHaVccawQ0KPaicXt104EPuS2ajbb5dVNfzw05DE1pjYqirUIwY5qBKF
fcdf82vMLQLObPhgiMDrtJp73fTI7Gm/LBbg+E0ztng9vUHmWd+pnBtLQR6A31rjm+xGe2nd3lLp
nXILDsNQjCRibEbYwpVTBuQJswI0hJcBCLBe0DYtLr70fUU++gCnV5Jx11T+3zSAGbAwq27RBL4Y
hp5S1e4Wj7Ug03mICSXOvCvRwYea5LWL8614V8mpixp9x1pYuPlPQDl11mkMmN2udSPm7etHjW9p
Xfymg/Yg24FEp4antEkPyhmjoXaDBnlObL2qgM/VCrtNQ1LDJxuxv6MwzX8Q+hzm82h91KTmBRaU
fDOOujkfpKv6rI4tngWdLmLW5Q/uGXCRPvoNyGxjz4qmcrBoN3Qm0CcU7MNAQnI6967/f8EG6Vcy
snWIZNVcUeEr4T6+zQL6tnzUGDlC/+6O1bFnbWfn4UZRZsz+PF+mcUj4/S7QMQxiQJFctULA3MM7
BW6uImSiDwmAPdtJminStkp7iMclr+abIM3Mi/t36I6CU3eMCfhZ3QGOpyPbQF+L2TZ4L5GdVZTW
3BxXoBObTflJF2/FYn0afMk6E7qieo7IJKxJLd2tmAGGH4GGH2p6tQshLKIV7yoJIDhUnr0W3krh
/VbkIFIj3f8LwMEz7NoJtwSM7LCR3ITOsvYWrrb64syCiCRmrh/Q6unCdnJFoTXubCDzQUHbhehP
g+HDruACMIUUo8RQrKkR71dBgiAusv9xkf3/DDpGh4sTKU32JEBcdKecVS46pCNb+/6U4kkEKPYS
cL1DZWi9xsBrbGMhXF7YzVeBFu7AKZXMuTzPEEM6CfkAh3OvX4G2lmYuE53jYyxO48pmJt0UfTG6
uIuN3z7OipI8a39vPgFdYSvfH7J8j5D9EPtw0LtGqvQW2oH403ryYPQVysT18xtsxmuqiVZT83Qv
Qxeiwc5H9XrUPr+XoAsVV5ey49K/kX3o4G9QEkRHrm3xEh8saKme0iUWMmjjHQhI4upOfirjybt7
Gnz8l5L3Q0Rs29g+Kp6FsOk8camqYqhdwhKdpQLOGCULeOkNHBn/UVzxkMgaVYbQO5ad1s94AzRV
6/R5gmPicdmJcvMK+p/H7qeWBnyGt43AWtqLGJ4FgbiaG8CPYAvGfZTzowpSq+SGQV4mwhplquDy
HYQHOURYDXDpxu9BSkAPa2qe32G9odxcAz8PEl+EeV9gaIBo0EdCSzJ1huGEUOvc4wyP/xDaV+t2
3Lu/cmxMs8iEvBtIBlanQa/nqIlNdKJYZjApK04H4filfYFPN6i8QlPa4UU6BrSIFtES9C4rjaVC
Dy1bTyb6tv8dSu+v8nJ8fX+bipaUFui/PgMQfR/FU6htWN3gOasEU84TOiQSnEIWvE0XC1Qj1aP0
h+c9+/8/L1cjGwTsSe9ENcWm7hFOsrZqgEkqT7kWEtGYcSZba9ciNHFuTHIjIbCfDniS6J0pxg4l
+SFqyUx867pyUrj5qxOXYRHWZMoVYwolyMf1V6vv7b0iegszvvkwR2O4VLBewUs0A0/P0EGZkJwg
/aG7Fh7hGJ8/TB6di7FtTn/bfyIvadVdq1Ku+HDp0EAYmuqSpZyOHHgXrF2bsnDVb69I75OY1J9E
v1bw0PMHXvkno7rkAy1p46BS4iGVqSoaVkmgbiHAY6vx7OLieiCCTZ+kBaevCs8oW9RChK6t3Xop
8p5ln7/ycLGLa19I7QRJUQfRLSFnXt70E3EUNyWhcE+hp6XxIURUrjVDB05N/a65kOZc53lRfz6R
u92rdjdOFypdMroSRAr2yZW/yQybxH/hovwOI/JD4gjN4VuF3OZzHaaYEC5Wmr0M4LLNZ+hOG8SV
nsCsvJU82RG57DPd3dERWmWYXqW0i9x/MPatdCg+kOWUQ6tD7kc4fOWPp3QIAPbAkUKxcXvPImJY
llB03FeZvfwQL5T2omwZTU/hWJ+drurrr1jdsGiF2HNMqUsvFdeDxWNsfY82HI1eTXiGp0SKRkoG
7UgN5PC8mgOK2RWt2r+cPmJFkM1rCncoPiDw3pBCjfdKc8Zg5ewls3w1Hfnn6IUUguBI4/lAOuVe
xD7asI7lC0WceUV4d+UgSVnURscLM67OtvRdDoEvcSFiWtzgWETorctigMkVBcUK2Hi0CRO3usiF
8M0DZ7fADegWwP5/ClBzLBY4ImIRJzQi9XLA1REnIyRkR9wTDwL5aR2zovg48zDYH7kN1yBCF6Om
FzXPD+WaBCgO7n0+5SNJBQn/s1tzgC0ZDJNdMhACUKJvtYuesMONmC6iCCPgxZS3BhFHyunjOvuS
H7RTlraYg0olZcr7buqbwSa6yNTEgYemXILY9jQ5yVYoE04UtoVY1r9+3/ozeP9nps8ZBlC7SYpv
NUpx3xHFtP4A7aOnN5Tl2QtxP+iDC00BlVmzwNZNFNZEERmRGHKC///cfZtsI/XF/8tSVyO3Dq+h
TGw/Iyhei7CeAduXc/eZTtCtF4lDSQ620U9koOJQm+ZbW+JPbFTwb2gM6ZIMHzK1I1MV7tCQ3vRv
hivDjxK25OkKFwdOkHebW4C0nrSW2lDUUXN6AWgpG+zXDMtVpfJ99GGoUVarJS+7K1aKoU/pNSO1
GPij2YS80oBWv5o3NlsX8BB2oZlDwGooafZFlKNZoYficvjV4r7BUdzYjxk0GH12LCWqIZJ0XA1R
smTP0VO0xrUprFxwmNDO6wqb0FS4qp8ts5oXUE9nO3U6aOQhfn75V+3c6NNGb5NwcRkCRnJZ4VJs
dgdJhd0wrJksBs8pGNGZ4a+sqoORkciKYgJAH1jfpwcCxJN3YutExm4Ptwhw/m1JJlhfHPLKxSbI
uoHppMJ9Q/EeOYbIfG29lJo+93qMilx4UsQjEnb0GlLvF838fhNP+Ahi2DKW4E3DxhPQ9Con5x4U
/ArmaYT73aCHTBqmB1L208DNKMPnXvAlLgw4q6/zQ77IoY9Fhmuv5WCPgCfMVs969VcAy1PEvLsq
m7A+wv/OpWMOMhMIVS0u958ZIdf8QIbqvLVVOJdEyDVDDPWuMDLfhKFkGW3WtTlZkwEbrAbfFyfX
c82U9WUxi0D2981pjbSoJ8sIWRzR8pqM473zG0NV6ieiVPQ3pvmH44RSFQM1/+Vk1fOZqOtmRR3+
nuKiJ+vXb4+GByS75X1HVpyx0I+CM46gwJ6RDpuHnCcDJhrXuzytqPj8kPbGn0ZGWqUalr76xGKe
lWu0cNPnquWHRUcfWZ/lBwdA3lSVl9oV9+RHCOvCG6v1wJ4y63v5KApz7Xa7U5VePUh/CbGKYjcG
scK7DaT4J00Onn483OeAAZn1DO86M4Me0m4Uz5uJ5bPShVykGuDGfP2yZVRlKClfKldaHA6S2Txh
pRbwKije8dcZg+ueLP6r9brilWAbSpm+hc/tbCyy9Cw7BDK3Bqy5hXq8nIBTaT2Ib4PzyeiFtIjV
9lYo9kwPzzUkeNonGbGhGxFFbP3GrXKYy1QeJKFxefU0BKb0CjrItZD7xtXm1B5MekXRwyv1v88u
/GFUmGHQryK57KcY4Fzbu9MTE5kyGSkR9jmxfQdWIPiRlyyQ2FynLoSeEbiPkzC2hT1D08SFqHi1
6Z9rr03vc8snkJtuOclAu3ihsC3U7vqE1aCdotoBGMORal8UPC2tP4u5RNNnfxlYaqIHpT/8OGkv
al1I8W03ah8yVNhIdj8tgr0Fju8WMgBlPatNkfpKqCdJwYrOmAwFq3jBRyFN2wJH07YqNXPETixd
zjD3Ki+fVgpRJ6zTqx3MHqA8LeX58+QrS79zUgSUERHzjjzRDIkOBwS21pcucXn4XJCJnxaZ3TEi
lvLHg+tLMsn2nLZg1Nx8nvMN62OPeSX09D8gCTGCyQv4Omiia0ZuY7biUH+E7mlDgo+/zrx3horp
8kTXVHftOLHW0SILn8Rh11AtmGb0VOjV1G4YAGfbaCj0hGKmRc055qs4UqcSd97VNRtL7Yj9CkFF
aSHPcSYgrN0odLYHgT9GGvWtC5lTvT0HRRVxTO+gP+PgURkIzaZslmSv0KpsBcR67AVB4Z9T1yRm
esZxW7GdDZ4HtugLxCQkbjvuJdT49F6WG3dZQUBwtfKznHmblRsltyaRhi7dhoncih2vrM5zunwo
NCwlIyxrDlDCKPdx3iW9a8wRF2/sLDYHwsgy2yPsYNxsuuNL723v6vTEW9TrnDi9QthAm2phiHxu
nT9tH+s+saCTZYv4tqU8WyeksnEVNf1qDMwbtx0eVHG0EYKNBXcnt7C++f45Lu8Dng6Jui00jpE8
R+CCC+WYDNPdun+sfAnqZbstc29l5cDRvgbG9Afr7LW6Ic4kh4TV7xcS5GyCU5Mkd2JBVUYD78eP
BEbCdJltNk/YItsuirnh7g0b3LJV3OWqiDQm5QcMfQJFNHjoM5/tV/zpiUT9QT0ZGb5q6yTVQb3c
hpiqSPGlwgg2HJ2h2FD7L63vQVs+0MIp9HvM9DcIjEK6e7r2V1E7V/YFXR6+ZU+UNd3xJ2pVXSfX
WlQtf8sXpTiOsQmzLN66+Eq3aj5Wq/g+zx/SL9w8DMy11xWCqx0D0RFCl/r+ae9Zs4S/sOigO4Tf
+0ztHUr1a55tbEyD56rb3HqyYmFH6DFxjgpzZkFNX7OSqu+XlL89dp/E7ywxxEBwU7iarmexKbqg
1EUUKIku1LhkuaIL69HfWcOtxoIBDiGGJpva2wSaRyDguZuJjwGVclAxNoIrSaJhDFYZyrxf484J
bOCE2+GgdMn4+9JbYCFK7cegVyvSgS9pTO7oMc8ML/MNK1SIZohDfZQ/aThGHO9lXlleGBMr1MNK
IMAk9DCULS2K0hm7XVn2x763q5ejlbbYIoFqlw7a04tsbeZN/X9NdbmZy8kGD2jAinj/w+Xw+jgL
QN0KjzoZlzXCfiMbdAJC2hgr5i/uVoUSzeZJR/3w+hPhOgXxwMk00FGxYa3iTFmtNiMVQkm11BIx
+Q3nqX4zzi6t1f0oD3Ilff/slU6WiHJkJdXMBMI2RLtent9P1HvSrolCv9xf0pkYP2IEks+9JBgl
W4B80GtWmvyHp1x1akpCXOFJhMGhoOpclfFuk6FA+SY6IbtnTMWidokgVuGqJquRD+jNTThepmQy
RwTJOWHqsYU3++ODjqOTLPfPEsl5loZ1vrBPAkjvbX5TZF0W6y/DCXa7fsFxS89zlSb1TqynNx7x
7pN2kHX2VEO1iJO6xRKjJ5E/z3cjCrayceszjB1dK/jikE7Jgj3F+ypkmJo9/MjuLbXQ+VeTDsQ3
/OIMzwizMNWbCp6cu7QwJD2HSn3L9wODtKPTG5/lbrJpZ8TEMaq4qzkmmhTpZN1GmFYSIofZs/I5
tfogpmAZZ2duSSnHEwucUzuhJHN8I2ha7izY3nmAso5pQ7gJgNKhEhjjnMW4hQEvsr5W6f8DQ4me
crHc2Iwy780tQ25Wj1H90Iu3+jsJcLfHAX6WiB24//q8WrKRYJLRzJFQ1AEaRfnXzTJsnaA+swIw
+1P2azCArMfX+tUKZhrCTfPXGfUZV1C5sz6dIEJp7gCcj2mrLuj+lDx8v6hYxUMx2lxWdkp0l9CH
fRUwfemzcF1CTZKDqiSlyiGHMwtgcvp7OB4H29Bj+pdilq95Cifc/xhVX5xAgZO6Dw/OxuIUlwQ7
tXl7IC8C6SLJiXFJU+h0DVooJwnSbhdBrzt2kjdNanWXzCzVE+vgt1PlEuep3U4biWHOySNmTl5R
+Sqwa+ObDlT1BcEJBS4JBHodP6x34ZHxBijq/FYq8YsgUnNlX70b6DmnR0elS+i+8/JguxlPk9FA
O0u3DE0rfN4qYWxy2GCC48qPgpQ1ayuYQuOB7V6oeYw60JOLxi10HdyE6tBLSSLkf70p4qJFvc3d
DSXIHnlEvNIgx9h03M7fmpBlK9FzjrpHsjGaLADtIMSS0ZrXRcUbp1HsLPdkI+jkHBcNd8stPE3R
4yxmCc/bWpBnixY+2f673rAut0p5QRevr7QV3TAnvAh+MfhiqtK3Ro8G6M9ehx7W4ZQIOen406r+
ncaeZy8220+PFGGe99VCKKQ/WxNbx3s4Oj/yZ0mX6FvUza/BybyIbb8pAEW7aorlH3ViDxe5erOL
lSCrDDLO/NqepKAYoRh3zE2hJtEIVk0+KDMYeOmeWL1aNLWA4CIPyjOK5ZIx1gb3uWrdetjF/pbT
7q/HWnTCtca0blqqo0meVdPoDyqRqS2GTAZ7R5H5O8VlZW5tRXW3uCYW0LRvxJHpGxijziU5yrpw
hRHS2c//1IlXv2Gu98EYKPd9eArohMEdFs4dpiII12rDN4v61sjTdaFCrEbk97J5hqpnvMxve7Zn
t2Fdi4UqCx/mwUldh/oDQlwzQLy86KPl/xpDBpUW/qvoXWszOaKnfhHqcTxJLgdgIlz4BEb3NpJn
o8ONk9dlNMbh140OIMhXmPXLBRA33GtrJxJVfjoYgVXkXFXvWz3S4HzgNfj2Z94PKLU0c5QZ2WDq
EbOeOjiUmPLHBQxp5D4oU3igW9qfLrcjLlSRzhRymsA9pmjoznFGSWHFtLMhhkgey8B6eNPHYhRc
122gy93NjrkQidJpAWehzdoG+xZGT1mFP1YdPrZpTimlgvWONnYyg2onv6JWLYgbd4d6HOqgBaG7
Uktxt41y+dNk1caI6IsHxivW2FxsoFuVa6MSKbBu8qKxbRD250LnNaLHNDKQIxkObMIFMoNW2K4W
QX+ImCdUn6477er0SO2i5PoO8b7oJTbrZ2t99uejrHToGgLEPQkrCRYXic9IxcbPWT7K6y8X+Qro
BwP/MW78oqsIQloaNDRN4lANcUstsUEISKbyW0Ri+tnQ3bEpOXzYZK3x9vCVAu6uYR1v0oMk3fSn
x3xRRa1hWS5zH0IQ+NF+g9G32rdVqzLIxS+P0czpWdPZ1MpmekiMYyUzOK9srLScj9LBYQcUjXPA
kgL0xO/csWSB7PioUBDXeuOc5LiAO1BOLpK8gPBIXuWPa9dVStMt55OZR2SmZxtCdPEq0BQzIyyi
kuKq2vhJfShRi9fE2/0iQcdfS5dIdZs/MbyXWbhU05kWrVMEOCKtuaiVBLd7sY/T11/OzvR7sD/3
B/o8o0jua4zVFtrv6KXqQhLtHfQOlmNl2Ht20TpsSR2DGHb7f5rHVV3Yp2rI8mSuXGupZ3p20M+g
6/RbNhtwmnZd7TOjXJF5ya9aaQJqcYbFhI5GhiPsm4zb6xsfHSgXQ3zpaLQyo/tNLNyCe1Fn+z0s
J/ak5u0AQeGLhdNOdXsEnYQV/PG9YBf/ZOl/rPDN4b0P3metpyI2eCSj/He8ZnMrYZcZtxKGd/8h
nb2qLRYVTlYLp0GxFkFUMNNjDG3UmbMq3rpSrIXy4nPMQJejxjNjxKPWhdyfJq6lEifCM6mXSYzc
Nk/8GeSEuDte5mvuieIVdyzLgNAHRYDZ/kraXQCvFKzUtml2BNOPhU0OKUTdv6ZVNEKsF9wLcJML
koLXh5e0GEYXrDMH0PDC1V/cSEr1bWF0PwWWzVmwR9PostwTIKQSlyfUZP2AFlLK79ItpMoWRqLH
GAO9xQ5PK+ldLG8FPOPgNc8gPS/BosWozCynjxcdZjBEObdnyqS/fQHds9Nj3fxDj44PvkN0z+Ea
8NWBCVpy2rY+FVwC2N3XBflTHTHwgYA5XhAW7FXXt1a9We95JhnzGHODJZ/lL6jekR21rRp/vbIY
lWPbpKANYw4aEg/ToReZLutHjrTJHqF5SfK6m8UZmLZ1yMrIGVmB4u+pEI9FPrLPLR7AjAf25QXJ
Lpz4dDCOEUjONfOZswX6FFVpMxCe0IhmLsSJagXpXFKXbVh3jdOwPTVPOCE4yVTuJPtXm5Qa3e+7
qjjxlP5j4fK4Ze0S6bq9YU6hZ/JV1aejUX3nuem0VIaRDSVvKbueZC9nzaCiMkhltzWyDq0vtQyp
n3F7mJ5nMD3Thsyiu3u4v4cZ95TFNaJ1k4AorGkWOMfWlZ6nfEAcPm5YTEFkVd8mjopmybyDWUwX
nc5Pj8ZlTIF4e3Rn+AaH/ePfmaWcAGydry/24QHZht9beIgbg1l4nOZIAm/4sPwbtMSrCcMrhP6X
9YyuaD54Y1bFZtMq8qEnfE5WgsD8ak9RG3kBTCrJsbp1TsoTQ+s906XisM3EsZSfl7R3hwjN4I+N
u1K2L6NdiJwgKz5x0oykHGIx2Z06BV93cMlxNjlNd52JBTFIqLC/bTr090w/1PC1LPqP/f2l6Wrb
vMd2TGVziwaW2RjhO8Y1hsbupSaPJwtkOJ4ZsL3Ddc92oQAmjoSJnDjClZhQ+PYEcl4PGNrH+Vs9
Vq8w2YXKLfOAsWdjjtt+u71gFvso138SZyaYelWGS/dtGQaArYssL66+vLVorO9OPz+NPWjW9KoS
9zL6oHUlpj3+zKkBCgGUlFQ2NxGFcejVBl+d9/IQAREfxxhDvcKFQ1b6pZXkEhXxs/feAv3AcZzf
bzIJezN8rXIcwlQNfrq+noMO8xi3EWLgnk5l9MuLVTh1PoYpb8+9QcwHtXFEXBmrsai3xvlYGx6Q
MV+a+eOppJwtgGaTc6kzAyrWEIn16X/LrgNhbSCyJFlnhnVAsdNWfSqkcn0vltIMR036FAqrtyih
LVhxewNAiejIoAWsidjXJfRLJHqj8NGwR+rwP/lFUKnN/GTdSjT8gE6tGB6HsaIndh7laZ+x9trl
nzvqmTLBTt3tIrDvJYhkWtiS+s784S1rwRDPnLpvubpSYfbquGZBublHUx8tMj5jzvCNvDUaiDKh
JinzGoThT8bHFPWffHj/S+2zEJWVU8RL5gyUPLjbv4UArm8C3E5O1k4/6a5yUT9pIGsfWRvXCzh5
NERa4gMzV0MfyQ+kQdV4+qneb7yKI3w2nE/vELUVPZoZNwNVCxFO7p72b+qQwiGjPEC09ZglQO+k
d77RBStNdhchIyuVmOfSJdY71snk7S72Hg2xi7Oh8sKibnSJmvRlxAQWH4AsHkbL0LZbxPHj9mN5
EYj8vyAlIzBN+8E7jS5hfyCivi0WMiOHhw1z9faiOLE13tKUckiiXr485IXMGQiLL3IyOo9T9ZTl
kdeQVpNHlsdhyI8CqiwL+5Xdn3maaLdLyPw4Sm/OZmA7KXY7u8er3ij6smAdyIPUyjndNHG+F/cB
ey5TunlsUK6KS1KBJNriCbr7FPVWEodMk50aasz/pc07SwMNZE4Wct6Epc3r6MxXuX7r1aIXTIEi
XnsQvCNvh+AaVE2Oz7o7B1vO76EAqUpMTWdVRMXryLhn9+80RbyOm9QmYZcSUohLSYw46sMP3sFW
z//Vc9lRwfqKafBzpUhbiMoqeRDMReKQyv1t5V2IcTWa9bd6rNK4H+CeL+off6PhxP7CY+89qShj
p7E1FQ4iVs3/HDhgoZVbYv2xfSJG+Fy6IilJuLus6MHAqHKGHVLMmwGJz6i5X9NeLSvWGgROBrTM
FIBCXy5dyTF3ZUEbfYGFauDEg4l+DCKZhfCRImYlXxAqsdt9scMKk+nKTe6THJPA8duZGPFR8jta
nmro+5k/dZ9ODKmoCpITwaime56HjC3U6lln1oxwKlDFMXcuTGQk/wj7wo1oBJ1eVmrV/dCsoLCw
+6wlJsf8RqwZ9oIMQgjffLsaY5TiA3XKIRKG9Q3o9hx0iwa4kaLgTWhIz5gYjdmIvaH+VdFq0sPy
IweBdPufOI3kZon5IiUC2H2K6uW8ABILTUEQS3FgL6Q6SIOl4CsRz8PoJ3RloKfVI3jhJ/t1BKVx
BpSjquiEj+l/xmsQkU2/aF7/tBO0aYn8MOflhBq/VuKSI5pFCMHS3eJzASUfDXwCU/4+0otuXuxc
3gdilRe2FH7gE2llqNqGeocEeT4mQIj1bQZLmnaRCnJUayFAOL3Qf1JtxTzLsRlL2+AomePma2nN
Id2W5SxBglDfQHxMcjJrabr1+0rSPu4aUEEulENDs9+8D/jwQ3jJBBq/n4FjmwqUvlWNVYn0w4A1
UR7g9wlZssafhIqckEMcBUs643p1gjqFcV75UjKJaLrgZ2rWKJ5HgoYSD+aTkUNsWqfEfO9AnbrE
7IKnM5cxrgU2am67Y7M2k23g8shfEIvMwL78jHl4hEuXdgVVv5QMYWEUMuSAtnKurNyAGxuHqxIe
XaYb6CToL3e2SGtprx++QguBJfJl5BkE9ULf2aFHbKrD2fpUhqjdKNdiq/UNHQwoK5bvtNu0jqta
owcBs4/rGlaIqQcx+yCCeRUoHu6FdFWo3kTfWZZ0B0AtGSev45qZFmPdISIqMw5JdtTonS5QTbdq
R4ryXwMMpIDInjl08aceTAoN16oJIGbBiyNniXwA7SbBfqQmi7Zh55nlS/czwmJh1Z4Ep31+BBZc
J5WR/LxEDvTrVN+cbiCcG4hd+i4rkX9+KpUD5anCWCZsy3BYKFaeizSfGVMtVklsooSQ5xJtrZX2
T76tNzT0gySWaQIrURkTNMLLodfJYikcBFmGw5cU9HU2TlbJzE6RfBGItRLGG2QZTDh8rxihbGW6
WmTjSDvcV8A4LuWIzUN7ScBYw8JT+laIyLRWGa6ViNa6tl97q7kZIB0Ysgv2IeDF99C+2MqiHjJb
TKz/bpe1RYRYxhmXV1h1Oit6/9Ny/EkTzrLoYspJ5rWiuC9ELGrr3M1wqVrqr/xgNnW73rk23O4b
3usxKvIdQQZ/54KXpyOXfM76yX10MlUicu+cXDECENN85zlDwRA0D8h2gu8+18WoAS7MtxGIResz
Ze96xz9kd+epmu8Ucf/EJSDwFxu0Q2ucgzgk8ptW/P25m1c2RLbPNaERzrurAUNBCiu35eWk2Tx3
A79Y6/a6AC04hTHu5gfeOWer00mhorTDD64Z5SxVKXX2T2Pp98gpUR6pdVREmEIA/9mCVdXRpCLL
qSJh13BvTdSvuXvDD10iEZnNsWLXla2ipS6astPgOqrVBU1MsCGrjxi0XvTofTH8MNsk49g/hstY
gE8KmUW+gCVWc+nAF4ub5nkGwEWBrQD8DnaS+ymwP2g8xi4hzHWU9XmFT94sKBhnRlnACwJjTRBH
4JrFC5sw1EXILkFmCznUZfKpxWU//uSDfjttiWO9SRpf1PSI90+LrJcjycEiEgLaPrsLU3/fuD0i
ksNLnDtA+7yulGspQdbCjqMwF7UbsxXLUTLRCgcKnnA6pYjfMC7iDBHAb9GVrHlNNOOuqfKS3l/E
abZKQcM4V7CHy3h8Cr04gWGSThUr7XH5WjsBS2mYfJMRDvtjclQF1bC/0WyVD/nl3A45u/U1pj8R
FNAtBLaSVdQgVv5OasNN/+3ccQjP8qV9TTCrhcXsCtJrSP/TW0xY1pQotaZHXn6YqH4nvzkdiF0c
AmO0Da2JgeQFXa4liVcn1oswmKcdI1EzRhh1JMbRY9waTLpxmcgv/cLXD2XGYSoc3fo5Wkwfdfkz
np7VAS2/HwpkU4T1YvW6KfBaZ3yTcQ04CzaVFkivDeaWCDACiUOlahS/wQdFzEWc0NtEqaJfkbWt
7B2I4G7KAAM125spZFT28qmBugAYzs7v8U3SvTUa1IQqoU0gy+X1uuwl+qKXuG3JVaKWO/2kcIak
6uXhpznNVrAKu+rsaKQ4MaMaCw5SA4rIUltAvzVTn6/iqujGEjq+Zx9vD/8v/D8SfixzLayWVS36
sais5EjtuUEd+k0dkKV20NyFulPG2bDHOsbz1g2Sq9AzmlV3/b7ojsIiVW0nVvDOTQPKYwvKUIX/
natnNiwXE1/unP5DRKmGSR87o4g9cjBMsN9lTvc1QYIMHk/wu+IP0wWWKYhM9DCsFVaKUrpwjRpj
D6H6M2R2efapoSk5iI/+OuRLwmzLalt+tZgxi+qGbZF4CXZs+KW0tvK/zYdm7SGM4W3CVB567hAq
/BbwuXZl45sM8dD/XSAWEeXAqQCsg2Pc50KHnU6WFw03DQs6+46pR5hxf8Y2Ud57dQvKZlQa+xOq
ntHLcSpSPnA1Rm0bkSo2LZsZqE+SdPWFmkuKyyPsC9MK2lR+qg6myMDlF0LFgiFAd9npkEGfeHTP
mPhy8p45Ubdsm+VS3/pkaNqE4XChwNaVKjE3gM5ndItq4gzyrjkkdB+nJoyVbzeqXI9OOciCOjgQ
UpsGp0ukG8iBO16MQVOG9hE4oJWPXvtVgtClXInsSI4CKIer79y3hfuQYmBsDv23lLjdRiHKcTyo
bayuQYx++x/EgBFJRChFBcUykVwnRZ38AyrrhlLtf9w9SPM8lAB0pg+224Ad/Sj4bw3H/kzdr2Av
t2sBaEuIxyhqW3Ad3PMdM5Yi7sGPkZ6lEzlRzXxYRLU8rmHHj2X6xmR0IIU9eHGRKsNORwM81Ja+
9FI8FSs0PiZ8JE4nDipVxvt1gArppstghER7M8orj8v/xjX2lzi1g6Zyev0VeH9QdaKfyX/6KJcf
hyL9j57PoVFH5mbriTqkwgNp27Fspa00/MEV/gdjNX8lwaqHb+xIDqpOnpWxmsfxV7RlsCtZ4Fjs
e5DohM/b2dsP8ihLhQsBXsjZ7YRUVyPV6WPA9wJfhYNfYFZ3xpUlmQaOUYWQZy00gBBw36eyac75
fSXx8oqxMw4vIFK+Ix8hUZbZRwZNc48OuolM5zYfblNMJSzIm4cUxlwRKKkETPt+a9JP2GrpQmdZ
PqrCGEBK9EPQBdwX/XdKsg2PWx2eS8e1LlF1Lm+bzoZU0ipKSo3nK1Zg65Ppsemml2/G89Cw7ffF
zD2fXtGD7qArFhKr25QvZeIf2+5dc7IrmXmsD8VNcJY0JEIpsoKM4gUF14eTD8SardehCfKWjvYi
x2+urud9NQ5khqJFrVDUOX39Cj4vxsX+lqx32h0I4OWJe4AhJ5gtLjdhQ24ZnzytUrj1tBWoVu5S
sC9hPup9GvFjoJix35lPjea1PwBi0f6Ki2dJoJ974L35Abd6cy4xgIL8N6iaNRoos5hL9i3avj2I
xSWlwtcy5p+t6CqD1+y1c3imywQel7evcKwTJZw3Y5vxUmOVhgokk3ZnUI8bURyh0qsBdlwGaLVw
+nWefDmFXuP9crCwaYN67a+RvDBsq3ni4FuYFW/T64KK0mKgcVZ4CyKeP1DgtML8tovybjkmEaUu
ZeRgj1iq2EMxZMqa0YgqHm5m8RAIFZIMM3Wqz1Ekc0LVomfJ83W7KFnnEsCdw56roIO7coCotgk3
HfdBShZNSBSonqYW7sf6Q9lSoQ3xn+O8EZyHOu0tJXcUnlICybQ3Gepnr5ozVtEvnFZyk9bTpHmm
xpajhPtCvkIuDIqPI/ht8IJZ0emwjWkZW27jA0uktCFhOvazhMQgwfUM9dn1qti2/8dChVWoK2EJ
hIOgU/9EJfx7KEfkpX2OKGY1AUR+t19y9l0bRzftJKucH1pOZ5+f6HDLZasS5YItgyepaaZpkcoO
LvqPUpzoah4lbEOmFqe0TDMIZRm9NP6XfG0LWTSC4eoIxEIuoIOqg4pA3srdhHyyW/oShIq4wpOt
RL2ZdxXeMwvmJBlocrw7xyEQ5zH6Tz+8MWSD460Tt4rYaW/5oDYgrDRynl7SFsGU+xvjONlGDncF
AGCXF+n/Fm4eH+FEYM8MTdsqpU+GYKWrDNj7R7NFNV1opGJsLa9RLaueI+mMlt2htY2MOujzOFe5
f2UaM3skY6JxNv3n4zf9C6Fk0M5dhHUL6HvTu61GLOUjOU/jLwbad5S9YtsmgMhM18l+qU7r9a2W
3l3XA8AKui4ut+FoTjwlcioS9DhxcLMQZ0Hkr/SM+WEgC6QF7mQiciQi/Uu5DFlWGnLQ3xOcNgd4
t22rMcBFToIxJD3WfqeOtSLoeRCuqHDJ9i5R1xIEm7pWN1cbvdrhkF0GkgARpFxBavt9BPx5oxyb
//dHIv4brokrstCCX8ulNGVt3bpl1R0Yl8Q9nAnW0Owkqbz6pW2Tdg+SH/GQXRBpWjJIrge7O7mn
sQAO9S1IJ9KBFZCu9Wk6M99wruzcNBtQVQ4dyEb04zhfVHUHnWVjY8L4L6k4BmUsjXvSrWYhIyZi
C3srkjEYhCm2LhoW865l6AR7sIJmDv/fo51/8MW7B+FCN+O+h+Qn0ZPiXlVKoTPZYPAYlqFckRbk
Zunx6Fvsv0oRbiVILCO9OcwwS+kzVCAShk4c6uXIGXJX4+Xfaw0TWVeZysWTxS1SE0U2Bud0SnX2
xO7lZA+WLIclVk1DxnSoyR3OQfc5R23eX9dhskTBlTct1uLkaiWhfF3D9nU1pnkWHDogrbxa2qwU
GmjZ4TMURq5LJnQVlf06ONeSGzI+u9PMrGQllMZWl+4FhgNTOeCDLjLU5mppp3vYHp6P4oFV7fee
DAiZeoGcivf6ndsZVywURuMGksXB91fPSDyKtqfIQe0gSeammLl68JGVoo0weveVm4uCI6HtxmCx
ZyEV3isFoxqzCKFKSrOHE42lxJ1BJn1bO/RYZOAgi51d5sVgNZUcZmcBo1shfx9p87nauUSAJw0e
OLhMiuufh2cQ0/ggNIFwR51cG0866YDE+95ACFU8fiaTKtw2TsVEyKzpXNqmd4XBuCBgWkX2gjfj
DE0XyEPxBagthwGpARas/XDzqCRMeF02C+P/p4i/2KSzV1alEnuF3LB7DD5de1xnkQNDPAdWFUkt
n/dpiefQeLpqauFb00kkBvijHN2bgDINZRt/kTiPPa+86ugZzc5GWBRyaDhoh0biL/keCFD7tYQx
jxRalchQQCOzffFN9vBnISTDMpqjWfjd3yW9Poy5un0vLUoHSMkEFLLbW0ZMisg6Eyls0eDBatV0
qo2Ly3PhHkkMdyvaooF9ccTRbCBr2XJF6wNAtzG0IhKThOQVyTxkXX+gWkiabJSmJOtuf62wx7e5
jE6Fh4DOVKvSjOy6ORD9pDSds2sNuDK6MDeztJDfHVZiYaRI94sT3dS/Us+b3Ls0OC+ivLVR8L7K
1amWNTQxtDgXS9BMgbZXYpt+DIyLOyMEgp1NbQ3ki58KxG4E4U77DwWTKHaGfJzaZlgpETDnwHTr
3UTQCTH3DcaNYle/c74JboG9ZdYx1SW/ZTAMOSp3ZrR6vXwvTIZjketjSlgGRjgDV4mtsLAeJoaA
v2QIJ4RLHZa6bVVB5vfje9mjbEOaiC8eo6yJJ0y7IYcnhs8/xCx334X9fGBZFdg0GCm/2bELNvxS
1OlgsEgoBZ1sAR8f3HIqXwF9KyNVOsd5p45gKEKf+AHgNpMoocf2YMlN1tUUcqut9vMh69qkkMJ6
H8rTz+kUvyq18gBbkN6kwbhbHDMclzH7Sjk/mLs7s4HaS8XKuNxxRmCRmYVvMRYAddPkMkre+fOZ
g6P3OLBQ3VjoSMkIIfvBvQAJapoBUn7jMF8BQVK+KiM6Oggnyp4k/grlcf0aeLdjxiGMPj9eRIwY
HjGSfahTHETwbw2QCDCX3+MEs6jlLo331BO28Y/k36gZw78/6xYIEU8tfalxmji/oBRJZsLTmwgm
2eEx/AYQ3Wp1cfv9SoEMBuV3ggnoAyILcRIFwzVz1Q+kjdWR1WxEtAFaiWAB2UxYdrvUYEBvsTcB
LoPVn3bvlJxQQvyZhO+yXYI5OCOkXM1SRCBv5tbV2/qyE6f/nboj3MTDaOrkfxljeGjkSXJHS5mN
v2QAgaD20VUK5RRMOsjTxT3waDFCY9R9q9VqLlAos3KI+tmJNhGpJMd8hHLDwEQzof8KAqW0T+YT
QFTby0Mz0zbmyfD03keYpSkUVX96UkXQDnL7QQu278kyr4J+e6mhGVyc0Nd+Q66pHWP0DzvGdb3G
MDADZaZw6O0DYeTiHqI26DCBS1RLQpeOLW/Leg7g7Wqk9KaeyyG0e27w3A6iOWyxttzshm1bvshI
8M0YwmDO/aygfFasXTM1weuk934r9E/zEZzZTaHSxWlBc7GaCCu2pHglwwWuGeTWABJ/30VDrP0N
RZJNEBB1KM4rlX/CsEGZljrF6oSqaHuwdKzWjA2MwBB67RbNK3aJQaZvc/JtcO1nyuZAmNJF4JM9
kwyaV1CHHA7UMwLaeQCtY1aN9c6EAQP0SScXzlbemHILaAa6p8TMVf+DSes4ytpjoBppwdIDqUqp
wGFQDHTUIMpbAgT8gHOiwG8V0XvYrvjQKRdzj/0rppbex+vhmpza/XKDCra0MZ+vgtirdZEaQHps
0VRQVm8Wv9VmDUVI81Ka3clRAr4Vz1x3ROTIYXKhWkpTR/rmaXAGdErCXJ93DbrNY5JjIewyyUyU
saQNmYAmewKtyN5F91DSb5ReA8ZYixiVqeuBTKqV8jkuvvKMDAs6CNc6iPdYGWiSrn6R/YAPpB8T
7s1L2e2NBpxrysmR8su+Odkyl1t7FfP09TQuce3ZrxXA/98licxAhesY7Gs5q1bN4eRiFiVuYRWk
13OdxATd77MJcdR7F5Ierdzzh++MVqBi4fwjl1eC8+qlLQeEZl+8kNsddHapITk5TP6XL2fS/qvg
ewVNleRPerYsIwHfpRsNIqSGmo+pNcLdLxkuFudJpCp6E+XySZl4d8XB4ftgkSGij9ODFj41sjFa
JmTnw67zc9GoQYZ5+iSd4zydJuRrIxnBkDx4qetP9WWBwoPIp7MS3aCCpQYpN+jeD/sdm7FxzQi1
Rm8SwfhMC5/RhOmcJiJZfqjvdGJWAfmfgEnSEW4vJh/IA39cP50gn7i0AnuJfyUzRElOQGc7OIrj
Msj0RFe67TsuOFHY2/PNWvmdOosyFdsS5ffBURPQxfGRtrWEl3If1VsphlVFu7nXa+E3Q7fzyqun
DgFIZa79THhZ0KRuQu22T8IyTHqRQrz5S1CpTiwjSXPU1zyCELYJamlMB81uZFX2P6opEVP9voL1
p0T7e+4KBYPOwcAT9R6tYkWTb186S0HHIsnwVDcoFIXnMb1jdZKawvVAPmxO1Dkt6768c4hIl3lp
zkWuG2s12A9XvBtdFw8ZZeWKH7NA8YM1uuPJKV6LSRieMSANtyw4hfMuStv+cljWAUJOh0pt3XFY
qKVsUVFRDMhPQ/VEdKPEL0QJT1RO6FESVt2N8xNlPr606MLlLs5ouoCKU2eeUnpt96G/xCG20xj6
65KTDWQUcvHxNNxGQyhIwETE3wetgpw/xwjlOVFEbm4Afrd9ryMB3JSHT8n7FQm+9IB/OcMwiaS0
s+BV6F26LmzryNg/Ivuv5+jGJhnbg0XsqQ5PDee98p0PYr6Qzpp/XzHA9142lhBMfmxBdm8b0n4t
7PF/crwPVZW9ImD963GtfP6Hbxla76nk6vLnFvB4VvrrTLmNrTo+57dhOfvGOT7Oe7ywMfq7shzL
synT+qubRM/tRx9BCTpsQ71KNrOizbxL31DLacg+XV8d6XI8Mi1W1c1gGhvNkA4tNZGN8MwNSVyl
NR/3rSnS80x+0Hj2KriODEsQYpYqerL+afxFBa7wKnkYhlblA6OgsRoEM6D8N3jWGHlotMPHBqR5
slH/+zOH0b//848QNbaighIgMVPENi60Tp+y56KXvPtrBN8c99abWaJpXeAuHKCAdWOvDPL/gfWU
F7fN3PTj2lQLCYqPV+wbl4RyjCE7hHcehq8fgjpGBGK7CUEZRumamv1favduUQPKxol6gozgQknO
gkbJCx/3h4B0RHrL4UNQ9ri0s75tFgVjUPR+LeV64irMn+4fEiN2kWqOPdu0epRRxgdnd71OSQWo
L+fKHsNFLLW/DB/rDbh52ZTrhAS7RrahL6HIsnjSeGtG/mt+Lns3YuvaDX4hs11FybyeOmyOHaFE
vZoPDWnZhXEDeKVRMwmInqulmIY0WfSoGLx8tybgsFF2Bm/Ll+7iTVf0h2clMS0QzSrgqqcq4R3U
chsjhvI6MIwmD7REsANP8iKb0TXAsLKxLflslE/OSQVrrtG+3SG1t9VjzODH234kQ4EoTn3PlKK0
3048ViPDtiKqluPwdhbs5G7m62Bo7U2kruub0BCA3iLx2DdgsoLy+9iuPuEV1oGqBa/JpOObL6R5
XndAyg4x7r5EGQBi3Wk/jGA0GECDEXR4I+HZPQtm8SkWxBLtxsv/TCHrJCVe0UF0iLGg0hjI+CMC
wQ+4Q2ZWebyJlVv1A3Tp9W08CpYrkoAyXdWK8zTUWyiQzQkGT+26PcWk6RxQJ2mR6cxUnlGqbBf1
5yi7u7ekVjQo/wTFaXNVkPBKXIeNWhfeu5ur38WSDoiVA3oDcYuquSn7gT9ngVVdtigWWkfhWd73
7+ZwZDFQ+aL+lfWq1wwi2QMglWfk38PHuHyggwcJtgw+8/VKfwj7spNX8QEo+QMcaP4HWoDuVixi
zoqcaraBmD20TB7Zy+JLAKABQjQhcjdIY75ITNyLRnz3skjIIkq1RvbnCjr8PcOKlxFRTEJqXBmy
wmjzNAZYYw27Vq+3p0vD6gXvHFqaYBOtBruqCWSIAysXVHuDR3+GNHRIc+7Rwkc4M4wcqqbwkh1r
DEqpv23mVXO7xL5ZeuQeD9g3Xbm4himP/nbIVl9W21k5AM1j5IUL0rrPo0ZCIFhc/Ruh87KeotSG
bhEAiWb1jhtzPzBRbm7SlCbBuS3c/a6gjTIx7zEhLuG497qAIiGI4wg9yap0LaR85/LyG8GXEjTq
gFXqlT9r5GS48ADX0F1hP3R4DrpJG50s/24pJFjgroTjgwzCTTPxvvzTCEson4HG5SDUA9C5J4sB
uxIiVLzvwV6hG3rnIhslIAih7S+nlwFsiav2ljlydMVeiGrD0ma+iSD8D29Caag97muUO6MnIKZQ
791zol7f1x/qbN/JUcLqPcJd0Ytg1p+kteIPqoxhO/WdTBJ6u1iwf9U5qqYfsxPD+aeh5JAQzZiy
imupeYqhVG9wBHkya65wxamHhRL9/qhf5mDe9zf7RWZu8wTBQX9tJq48/qBTQC7wO7RyKMr7tMdL
FC45mkD7vNInXPqX8AI4ZYPlmaEkn+a+R/CHE7IDxNDf3bD/humTzvbvS2S5HI6ChplS24zyJW05
hoWJMDdRSkyb7Cu6YcUcnJHH+UKzzFDlMFhAQBlMW55t2xhBfd+BuZ1yba+XSr6UzV0vRlFR4PTf
t5uvbaMPCYQs37a9pq+BcRr3UTus1+rHShqS6TcaTT59hVzF3AUT0HiT5a38STRqTIxpy2MqTdoY
W2liksTpCAUpsWvOEh5DxqA2B+eLVBMbLkRr9bRhh5YSyzelsjT6JOfNmYgmh9aCuL8NFRbCzPNV
TGLB27QYdlWsmqAR0HQ3CBoswaE8S+yCw4bJlKROWLb/V8ZzGvoBew+CdcoF7h+ndwUPTLZL+rMP
qIkiR79oOGUsPhtoutdU2p5uQq5cMStnFDiac6o+bl12m9q4a33A5+eQ/tCzvHdWBG5qJi5VKlW2
ASccC0cqHLfo0MQySSH4PhGUwnWX+AP+iDcG+wcHB3T2ENUIDgZz0+kb0BmlN+qTUStAvGjeD/D6
/Uc17VOTkAjEeZ7GQdAnVoFl/IqZNuk1LLhIpOSqW3Ere+T4CY4F0gRyUJM1sbLx7kSg7tM1J6T6
1L6CSJtY6ZfI/JMtUqrrk8NJwnGA6/hs7ZHzaFnQ0zPXMczJpd1Zwy85Uy4rwyN2yXxbtbSXDLE9
bUfhzZ3hk4jECUsL9lk0nfuJKYffi8y+Q3I1kqapoLr17LZcAKErpzb3QIGeD5SK5he4Lg/CiO3Q
NY1JsaSSwlUV6V10XsovXR16bB/Vzg6bk8Zb+xcEnZFTkf6nN8fauGkgaIdJhHMADkFQGA74s2yD
jFSDlZLKAcgY3GWLBk51A2CyF3u2YE4igfA6WqQnlfBCKT/MUKLnd1yJDuu+zGj/oME90Mb8CrWs
1z+0wle9kA6gcek8BsAP7OfOxp0Wagm5zILuYyyCmYNx1XutEI9jp4eISDv07W8hLNomK/nS6crt
fkLuZahsXmlvV5XJ9cNnrZ8CZHKlaFm6T59n9xPX6a7fN9DDnJMIe2KECkeYVJmYx4QxR2HNC3VY
rj3oRHlTQnrq1lZeeqOYZUD+x3vxov/kEHarSxXVr30bj3sXdUfjLyDozNjbhNxVv56Nc4fkQwYJ
V8C7sFLOKVErKwnHGng17wgvFLy6GM333ungsnjMvj4ueQVGgNmCdm/bM6ZBfMazxF8UlUwTe2nX
PWy83bFL0YmWFgdpTviBKpdORu/BPLoEQniYI4b7BapdG8I3Q81lre1WCtPzbyL5ty4jSftUbCqD
cKkLLn3WieWOqEjufW3opvDRwOHROaTRWVSa7ydvByIRuNcLOUUICGkNhCn/pflC/TIxEDdsD8bN
aqquCXVpZ6TRi5JQZcVzF5HKeDUdh+2ZiiUzC9IT8UO9tUUnVWuONM8fXo9fUZpuJefuqnpM1+0s
qjXUXa91yxExWh0/UmDH8J3fri9XHnaEcjr0qMPVODs5Zn/DfvZxqllO0l3BvIttPhL4lKu93PuG
7j0PNrqz4Rr18ByBRtlF7HBweqQtVpbW/JSoI4zdDO3I/9ec8X9eTyY/Ym/KQjIdfJcAPiIH8Vvz
c7FjHP2Lt9O1J3g8z/PU36NSLcwLyB3oz6XAXl/AKKpQURGlQ6BKCBO36CJwBho5LRbF2wMjP2ox
DdUyQW8nwZFh70kdbHGXeDaJazPIyTMNVJ8f+S/sd/RpAJIVYBwornBenDJbeb2WgzmyOEBx9nRb
jXu4zWMzx7RbpT7ZwgrUHm863FUwVAU6QNJEOtHuAw/XoO+2FiTfa1sAeRwjev34x36esf23euOS
g8mElAS1amMFB9Z9Z5LuT6BP4EwMCJUGtyHOntWCoTO03cIIZx/vfcP5HTYlPztn5Pgz8vPVXKde
LsHHphsKZTCUpPaaUqbCZebdFb84+4FjG5Gfz6eb0/xsm1mSEgVbrOk2yxTPDUFBJRJc1W2aHoSE
lF+zILIggj+Yln73nNK32rYw+FMiHKD9hWt3gMUDEh5crShWD0TcXMYrwevPN17qSDnJ6uF4P/0o
ZjCoz8mQ8wku5EXB2lR4r3aey1y7M2IzvZno5YXN0k5alOQ5S05L8N605nu2VpHUgerZv7niFjMj
S0VAh1YsHmz+IBbcmPbWamm1mVQZYhv9Pv6rQu1Axd9GqDikPuDEauLYNkQmt3yHbCMS7A+mGaCF
oqkf5L8Ica+OXObHhwntUj0sdlxZ3C7npN+L2GQPujd5Gz877IPsoiJUPD4RLdVLH8JpVg3Sm9k2
CuSRCZL5dmTYQH1IUmL33Em6FpLYNABFRUJ4UCHAz/TpwkgHMg4VNGne2Ab+wMZHXnVKkBOySbhy
mZqhu1bEQdh3h/k/ydxg0qklOQzoBww0wDn5i7ce6KurKUBCK3DOptQ7ReaDNFTM5wrPRIWn2KWF
Gr9S/HHHWmX3jfQLt3/auR6E6PmwbfgteXpGZs8XJsPmSLYQRZwAZ8FR8JsLGpPBhKhenonyxZH/
qF7QPF6z4j3Nh0mKFVCoitkIS6lMkwEb5Z1km5cDbe8Kb5zimF+8Sh8ZFIGPR4/bGV/Pev+xSXQg
AB2bqc/J8tMGvlCT0CIvUL5blX+11h3AUR1ifHnY2kMi2aTpBiztlZfozLXc42kMAYpm5CROd/M6
8RMIUDfDlEsZfDDYu+k0WKQ/Pbxm5wRnwPx0WTvzzQ60kzmSTtmLc1HzBv/0pFE4xy71HRSDuWvg
sGugbp3SYEfsbm1tMb/06Fz3+NpGPlUReOY4lSeiJYOhW+Ih2nLTKSCh/qmBRMB0fbhrTMX6CHOe
UI4rV5P7Ks9dSpy5lSj0SSMY3qXujFGpsm9ds7HiS02TQ7Xw+fyRf/v73tOFl2Vz4FnP7BY28lYL
wqS0lWiXcxvS5AUk2tYZkqCHD7I8NJ334rGfIn9DTyjY9ODxvh2NqkCUX3MAObMe09f0tbgiGlUO
Vo5ET/ze1/kg0gK6kiMGttTBZzKhHujbuImsPoxXTclKu2VoUXsl1hLfn4yBg5mH7uf6IO5/GbzS
HDILZJNlL/j3qFM/Y4R0B3dHhvTyA7bamTG01b9FtxAV3dq/RY7+jAKzr86tO7Cy0o/28PD0JGDK
50NtniW34B5xMzHWBnaF3poaA7OdGsXTtucyISOv87muX4CiF1YSTlt/xTmptSGt6lJXWgqIXmHV
qDpZmYqC4ChL4KgQi92sQKMvm3SsK8aWTT4NUpjJYtKi07iUMrIP0EN69/Ii15zzNopKwQCx64bE
z3ySUKK72m5mPKfP3UJ2YZhHSN1zbSB8ND+Q6yJZQqjbIs5uJ4XjPMtJGyUwzcbN545IfPMyOVZY
PueITrqV2eb1c92tjOLJtW3kbMChmNoQcdaLLCFyZxsDTvVo4higx6u5FT+JVmTH8FWDJTpc74CJ
p8qar4Ke1VNOqFbiTpsO78OoZgOuzvv/xdnIjgw7hB93uMtgAMSOKpLoUYZL1n6XXmPzdTmwUx9N
8gUlBeP2i8JlhN4nbctgSKo5WEg5IDzBV/X7IO+Gwx3BDe5iNNTN1PNAu1a2pwJO34PdnelKHDCm
rx5M4Mb85as13naHzz+iNuuD433PjY6mRiGXthwv40M9sGL+gdGid7BNGNi9xG+I87d7ZsCkjf35
CabY8DVZaD5Wj3Rjuk2XquGV5VoJhqeg6QGGvrWBkigEO1kqLtQbUbJwf+zDRS06fox9qWhuyItF
XJNBO6EfynakWxFLYUpkde+rF8roAkejSFgkRLaqxdDWbVzgM8IUYtqZWe+OpQo/SMpJMI6JFbmy
/WOPbMVoDkeAKSUV4EFbepDLIhoFN3uc/ZXK8gqem48be+it6/VbXYWgdhzwPaURzWm2z9A7yXke
9anip/SP+0W29rf5HZYXS3IZU1J1pJbvM/mn4IT1K0cDtBXL9wqu6QCEfPXgYacaRnR11tg9asSU
IKPm8Zj/0wQbUxlvZScK7t6h5uY2f9PYQGbKS0EO6wMesvWlR/Wh+Gqej/xKtaqZRY69WfdEj5eF
cLb7WvoymjZfng1lBne/1hCLDxwCymAP1ns4YF27/QUPbY9DrDYd91W1Gk9b4g5zYlKKI7xPFKJl
mTBMR5PX84yTxSltbmytvGF3g+TLLyHxGgLmCmwrUvxWMNEjjCP07H1yA1JkdZB3jDVh3nzAWhH2
4NkSUX9IVQopDQkC0V7kmpVaPCYL0lZzcB9Ibp9tLN/lGLCsqQvS3nGZGWzRbGFNyItWgZNMwu7B
k57i8wcPtRZ5DEIwC5Qj60V8boFMg9/d8K211bK/JkVUt9oBxw8CI48hUeFYqBJvInHgUjSmwSxD
GilRioW+oeu9rnaELXTuKJAzOhGRhb91x9kHRTrXm34bSyTidZkbWgEqvrfFmRaSX9alMkn4V7eh
MP3GBqJzYFkd7VHSihy++rPREcowSgnxTLKyPV0vRQy1Z74cy8K1MfFmvlRoV4j1r+TfBJ0k3Bbj
rSzmFBxFQJVdicGHG6/c4nIGRgJY7l0tmoZFlFiruj3nwyjnjMLjBXMDRFd6An5SvrrEDDNNBUxX
yUeFUZCI5O0QrivfM98g6H0dAN0Hy48S/GpmlFb4Bd/jl+o9aDFoy8Nwzlc75NCS9Aul0XBbQfHf
lQKBBxBQ6O2yXUaYFA4eSTNYtJnAqJRpi2qo5wle9IXDQ2y3SnMjEVwMv5vuB+JtlEtjer6JEXk4
BktTaLYzfe+TJHlJayBQf++QdBrLQ29t1qtT8GjERvOgNok/MPet+hjm1IqdMBKOOAnLj5akxo1P
/ZjsNKmWI6hcLGnzYNdPBgF5KZYe0Wy7AlW3UF0utCdBqBAp4vAtteRMk34ApxI4Jo6uyxStKOmT
tD1ishEzKlpnt+3Uv27ZjdT+Ds1HzfjwzNFQ3W1XYlK064BK/kIlEQKYXndXbErdQJKLKUtaRZ5e
BxXJBOKSIhf7BTXfiKTiBEMzwkNqkyRlJG39cLKD0mcsSHLp8lO3deKsgFEAiHPlZ92GPrlTBBIV
4SMe+h3et8KRTd3/iB6q41Rx5xedMGSGnJrfC02gseXP+cm7DXOvpy1/3nm1nCN/StqYkktEpncr
0WDM0k2OYA7osYJS6GYuA+95sU7K2BvU9i5pklL1etdSVEq5uzehTyCB9dShcOSht67ggcLjRrKD
uYU/N4LjyCYTjyUCRZ82rSkczGpuZVLSosvLjARMKHb8OE0S2oIkRKOMHHUm/GDM6TuzIWzWiXot
qpMdYrc4s7MYDi63SBAAgDy6hpzYKWF4Hoogw+RN7PDV11FCpGoHt9dOBJj0rW8A/BYhO4MHhP2T
1qhFgy0oER7UpAWqFstDHifX4e5BdGM3YKstYQHLlvSS4014n0ZNuVkchoFzGboB18ZiyzNxGFhm
Zix3dB7e802IYaBqX9dxCocl0vXAocce5R6Ze1ii0iplalCFm9m2d/CGTPDz02F/XNb2NJH7kkbY
/iEzDKqjsjanFR9ApYyH7tkwLyExtaQOskr5br3lOO1+Q9y/TxK6GzHS1UyM3dQt8et9hn8JhEDx
xqy10oVUHXuB/+wXRF28s9BsIcMEpvW00kFiLGaJ74iZHwIySwwY6Hi0JCfDYHilNS2ZCz8lWmvo
U4++8aAWvnjIJtsQolKmFjNQyxgTQq/1RLf5s/+2lQKCPmbvXmIeSUM8+8TubW75rFXrg7JwpdqE
ow0zk01R0k07l1CYPSKiuKSDlhnBqUMf6LxRFqQY9XOPBcV0tMHjplyrdPx5QGJgfnR2tDRUu5ZI
W/tfrf1HWQcFLZwXmgmWILPD5jWoEnkHnnDcQ5PEyXD03U8iScG4kcFdJ+FKAosrthAgTw2FZX3K
f9JJU/LHwvX5F/6vJb5v5pNwc++Vnu+Kr2kEq2M1WUX3jnzjKaSOtaCCcNA68/qyH1MPzkFnJMQH
d0PX7O4ozxw2zKFQyzVZJJUAG+dyDW7wwN+hpKSeCYt3ewI9Yr+unJu0hPChpVxBWDVGNKhOuptR
KIGVvCHkxYEtSonqZPqONgc6jfqKBObcbxyt3jnSEna1YNwY5iJgvD7pbKm5ha033fge6QPBB614
uiinjZzIcy/mQEOnIRJqpZqpVsFtsC5z/QPeEQh7S+F4r0v98X2NVrKVfy1DF2vnOSg+QkLCKdpk
HqzOwO6HwM3l8aSu4UBisEIHDx/13MfOTso7X1oXbb4wOQ+1fdsREtwAibZR5ZCzD+I/U+kp+y2o
PaxoLpiutmpOyGG3chENJhbZHwEq/JGyu8xzcfkO/+wq39KquDzXTQrkiv/xwidTMmkytbNYHx8U
dk6Fy8jCWzE7Odc1JC5RnsgSIelYCcDDva6LN5xiiWPm1FZT8sFzFZ2HgdnB0yv7X5a6sjNKoiL+
BMQSVA3mO9nTydxYiVppTlDjBefAns9gLy4CAm8Va4bnnLI5JzWbPX0ymMCP7tEKhTm2rwTB0oLm
crc2cLrX9PcFUi0PwyBFOCPDxDzOd2NGU03rHHlzVoM0bW6arS+fPshOTez0lggktRrqgfp4qD7q
F3DYqPFTlfZUARSoyuBL8R0F4mRAfZo4A4YS2Ushoh0hYRfZFA87nlsUrWdHoKbXFOvAkc+2Zsl4
tnzdpVMpG4PCcqCdhLh4cchrVMnpirGcyL7a7T6o2EpQBi4n0PpV8hOiuF4c3IWFWwNfA+IlRRmf
Zn0Nf/le/Ta3fvEkIal4VLda/rmT151iSzG+FjOreGK8hXdXNzSxdhWji7vd9mL6DKUHRRoVD6sr
WFKSpWrt6fF6TB4v2jKP/NlyC3K0mkICq+vKMPza7d/OPyCYflTDgukbpC8kJazF4vDY8/dZWkmW
fZIxbvFVl2uXy2tuA3P3KdVzej3OgukhCU/eY4Uuy+qrIGjhedsUHga0PGB/Eil+EC8S14b9xMSb
DrvpKgqN1pD72LUO5GBY+tB5f1PQrh/+hpSIMKGWEiks4ureljP4IhKQSg0A0L9XQgmCe3lOumMG
Ize1VYa559oKhzeWD9ZHii+hvfdLMKSK1hO1KXheNjTW4wnKJEenlu1T9cY58CWmGccxgw7vHKM7
sBsD4cAbt6t6iB3fD8iuM7LR3w04EQwt59usmdVvvVSylCGz3H1K5Khzx9tpqzDvlEIxmQgJgU6x
me4xQ7/UCRt0SFYEW5sgSVtAQOTur9J8bOHOKy/VsLuO+H8N9/0GD3cbFuUbsKNRDNZfosyaFQ1K
DDi78vCaU45f0VTPwEyuwm+BHlJe1AVhTDw9q2CwnkGn6XW0DDq8eCdgqLXwtoaGL7GW3e4ptru2
EdLVXsxonETZoJHE16DDkPcOsFCjqZzzIESVJvakh/7Qt/cKiVMJnjIXIqAK82tuMn0dbKG2NA3Z
DJYmJSX6JQQdRM6IKA9zJKoH0vboEokvhvAZE6VUkgy/3O9osW2H5JzEbIsgOuLLalYb+Vle5n07
ZtkNkNSNvCVWmfZcv9V7sTozQNsRGbPrYKdWhKvCbLHCTNMvqlQ75xnzmtm7ixEz/AFy9IYA1Gnt
e6dLM24RlFeLqoO7o+1TJXj9xN60eS1a0Ucs5IM0P9/ONeuLtkhZ95/f4AWVpbNg9KluE93DGKFc
fQ/fXrbvhHQ884RRrmyle6iM2/8QtjO+NVJDiaYj2ZJFQvNTVldR/WknYCYBBfW9sObRLV2wIFh4
AKSyimnKDQhO0Z2oRII3xgE7Xwea3jfUeQeEZ3ki6/0QwJu2un/q4SMAUFJhlxil8e/Qg2VLGeYm
ROshUKvau9Y59awbfwfXgiO0cFUntBzC0djmK69nwyUopXv2EfVaJTcQMqqUht0DZ5UOuwQl5iD5
gIwZXqG9XsuRnZC+Ki5bGJ1U6bvCT16Q4RgkmweDReQqIBbEI67X5U3Rs2eyYHe/qtU4KZp/C1AT
RKI6N0WCpencGmMFO70fRzs2fxZeCZunYXNza9gijie6A0Ga266Q1e4NOQ0OGx26haSzY5um7oux
j3bauuv1wOMC/rzySUdtk+GSI2FKrDvZR4XoyGHn+unlWRDpc+AaazT5LmRP220+X+EWXaU7atIl
OyCBxvoy8vx1BEOSHZf48Q/e5d9tBZF5jXEP569OdMTcI4Bp/VCxLAVYQjIXhD5gF+JH4UZp+9b5
1S1jHrlA0IxoV8LUlFlHQsyXF++aPXIY+HF9f6bXs5dyBgt92DBfFUFcg1ewxB3S3oQwlSExxxfb
YLHozmsZoIhKrFUA7gF4b3YpSpkO5SVCWUd/rq0Vs86xwbMIHs//mcKN67eOZWDN6dkoizG+XecP
2CO9GLdZLi80ph2RZb/YDu4hhfsV5pTwlwqEQhlaKDOTWRJSU/oIVJCZu2pe6kG9l6OAcSM9R97K
kqkIpL7tHJKkyXshbkSqKkkyxKT97aJdACYXaVif81LQoxwWWHouf5gz4ndYOsN21sNNxnwdhCU3
s+g56TaYI7ZaROIsB5Qtuwe0wWDeMlEivOXRJvTgKuvg3Goo+9XR7KfyraePU7x3zS8+BYpNf/R0
PDQu8cLb8MvXGIu5RWoVvWxCKlVMTeg/JitYNRXe60YxRL/ggsrPsSjon9lz5Fo9mA9FDXCdpUBN
8IpZTETrdxeFil4Y3AUUsz6unstxjXbBmGgWuWNXNnAs9vTJAvDnbNFE/uDCiIFLNc5ifUbhJsMp
Urd3uOK+3YVTdvj9kTlzQZNtcHnECbtJqeGbDEv4n/bSjejg8SpQsFI0z4+0XbjrsWvnIXUM76+u
xBQ7vHVsYoYw9TCo879vSplCZsxSKUNHzujOriFluZ1dywLEdtxogYNcN4pnVF2UzHBVuJYLFyjA
+LxDiZezrxnJ1xdM5RJtgczkxdDnYimGgjxAS/XklXyCwMYXXUKrQVFlY8hXYW4KxKyEIlymLJCK
udKbq9wSlLMu7gxKikS0pgxbADxFui81Uuy7ZFzsdmWddx9TonhiQ2qwZd5gtLuenednObBPvZHa
8YMolsZrUPAyu5bjc8bZG05xi10eSH7PLtSLdfn9SFMxOELoGEx6EsULRP2Duy6c9wOjyiHvEkKq
rtHkyBWc/1jtBiNv42SY32iYBjSiOkc4JmCr4MS80J90UP6hT92jEfMOfP8qdy3e6JhJ4NXVLJ8O
buJg9JJiGmREt6VDwT+oB3PFh/fg9FLJYo+G2f41BY6r2zLw0EEd5qc2kkmiCWrNkY9nyw4eRRFU
AVeX/jT6ZKjfpae6t4L/1VwTM6tYUnmtlfh2KyElRWuWgPhsfCcDHmZVRMYEW0U6s+v7+VBOASJA
kJbqdTJhow9SaFJigMAVuMljVPMxFpAkVCNUKqU6arYY4ah6a7x+01DbOYN7L5kjhYt7c2Fdk9l7
yCoZyPiqFQEl//cv+UrIPmS/IbmaG8U2VQz+C7XrhaQKMt669hQLdpIoyknVmpQ9H4cGbdJ2JuUz
8+rBF+BZPGAkSJNs74xysKKb2IHRoN8ITJvPKYzETupX/JnDU/JmGEPFKZdxHjVKl8/z8JtBiQL9
J+DahgK9jY5EkdomsGb4gYHTvWfm2WXWmH3ESsE3LRSLZlYtZR5yhZS9UFqhGu2fmYEqXw+70Uyy
brP9NZqG+TEUgzuYT4lHs9jwQhe0CxoT5X7ysL1cQOIAXVSIW+pk0DJTdsHxvi9c3AoboI58ZoJo
yRjwxYYoLKXPPqdHFRHnCW5NqhHJayry/UJ1fJnIbMQJ0dIt8a7KyKl5URYmCrk/VtXbhWyxFT4F
PYCYGMWExKs/h83AaNGUIoHZ9pExHYYiMcOaNqZc+etPv8Nc1ivIxxzHGiSrCbuuHbCmRUi+dxYN
ClSYO1T0NwQF2k86yPSMCau3JQNG+pQRpPKTvapHUz4HqUse9sl9P8knTLn0wGHAC0IoWEIDKg6y
04zDBGaa1xv8zyyuORIacjT8OyqKx0M/Yw0Ab6Ks3IjPzK1bMb1vV2RfSp0xu9CIpC30CwLF0Zgq
41E1cZTyr5ROHYPboE4pt2QpkmB1h+nTS26kv5Aae0BT/te+HpVTZP1ebZ3fr/gDsPaY/wHPu4oE
YO7GqeS91JE1A3/rim8qC+tY1UI9YE7WMAu+/OYug5mfb9FLYaCBDLW9nv5/fElBafowZzxPiCoE
1ISLRQNzMwu64OuCieTGdFU1gSOjJj4r+SwDLHN6fmwctH0NZpdEwJi1e2v8MqbJV9t70I5SDX6+
1PU82LXKbvgGWvptN2k8IpXZv45xgbavc5uA30v3rcIh+wQqetMTtg+hUSxy64PRe+HUo73J00Zy
0I0LAJcwr59Dm05qzCxryWalju2FNrASbuiEDp2rEhw8lTHIzCFHH5JoCCT4X2Zsh4LdvgpQYyTh
qIWdyrzHWFm9yxoHqMoQhAy+F3wS72MKOOZdZLRisWq/+492PkUQxfPUnr0n3CW0CMpoBQUZEsTl
kfkgigA0DxvJUtTw2darZ2FjqPIIm7JEusC9tUxcuxUakW913FeHUgZAT6p5l7xvL7e8iBFOOrq+
posktTsu5GAQepsG1C8wKwshK64HR9T4wysX6z5+15JkDMWlAiSXDLOtxAx7wdmx7kwWPGQ5jE7y
PdW+X+0Z1ag9OS7E2ENYAsmn1TCIbUYjcK2lrR82FPAPxcJGoYTc5R9o73et6kFAGyHEGifwfdoN
Kle5rpcAnDwdW57X5/jbTQ2PGZjRsIJ0gJt7dJkJZrWyuARB66XeJW4MgT9kjtYON2cjGcgqCyOS
VvRMOr6/kY9CdgRl8pJbvp4ewxFp2FuUV1rncpqqXxpxBzGBDQRcuRcQsSpRb0bZH9t6qop2KmNB
TgjRIebBOFKsYS+dQRn05tRenVirqVPGZFarBVdU964I2h2zfGeLD/engDaz86jU8E5dnvKO2yGU
zIHQ81eQ6esH4NRc0YrsMIqIKGIgDGe5pUBjIq3Jxs+oOBUb1nn4kIc7datpTg8fEl8BitlATyNA
ES+ofgnXEuGiB6wRSObBBnUCGOH2cUplncyo1y0b6CFbU/3rPfHw/8RghSpvCeHsA9HgCIB84fee
Dzj+nBIkrknaM1LyVOt/up8zNdhP1vGyGTtFGmB7DxU0nF4PEUpUs6hoB0BLVRXTFqPZ5FxPxPCm
6oGn5560GjnSm4VV9aIbCIQd8BRlZJJiS0Zkep5jJkpRmWO64Ed3V1kqOwzYb2CVfR+l64EDdxUz
VMLlSmJZ5v0WXg4tYLNu/P+AIxPJg5MJ/FUSRJCMSKO6PmdPlvHKb2q8F+/P32fQLOtgYWf/Vu61
43M0y7TjPw83xdQsNGPigZyKjmOEt5osU6S+weB0uCSJeJeNS2gFErpZBVdrOKHNnASca/fXbxmX
HAAtDkqfaskzYD38KHhZE9UrEM2dbWZBUox38WwTTxo7aH+qCBFgXTku0F3H14Q9278oEnoWFjTt
0d0R4TDTN++7tQwFXea0crchC1dtta95uO0E4gYFvEotdZGVV6X3DSkJnLbQk+SK1BYxNpxcMHd6
nI4QqGNpCYB6KdeyIjn0AfwIgdgS60xq6O5nvoIJLGAYIlp3h/Jx0kKqqD5L8IMQHg74EZ7RgctR
281x1bP+8tF+nGvNmBL+YoVXFFqhD6RmGBoquV0goSCLgVYbS8LJlFJDaRqFXqXKdRsPsgNju2Md
0kt1eMdIL68wSdKBKa7JloDhMoLUjVZ/M+NvD09JP1CaeiZYLoGnF34j5BUB3wxMjcy9E7UPZhN3
VHkPFO4zUDQqP5Uhzc63y99u83K22dzTrRiS/3GClDu1Uy5CsHCQQ92qLQW4Sj78r3wSq3mheoEk
UPQkrFaFSU0e8xME/s3fYTzYlhzN03uwZcJsiIT2yO61nfmLFQkUFnDsuS/sEiVfwyJGVdPKDghZ
KyGSx9pSFXkTQFf3MDTVvVtU1Y1bEoN4HDzTblcpLajC9zUIlKzx46xwtnhoFSTCnidyoN9Djjos
rS+9K1+jNkFAY79y3Wcc8DCv+5r6spdTw0pxSsHbEAC1murJozXlgtyvj+LihOwrtUBOkDl2LvO2
a11Vwtp8NlPvr2QznFU7je7Yw7lVkXqryzztxTmXtULmhILD2paPlvvrlKrqia6BMmgTgxNO64E7
It/bQRwCABOs0k15tTm/9pyc8PxKQ4S1hwYEHkF9r1R4H0cvCYK0zdI3J9rmrpJDo5M5QesNTWcA
dC8S6y3LVG5pTpaseEM+SBTqV1gCd82Z6PsSeEoiQHFD4B8asQdALA3X28SlKNhnr8i5mTia8U/h
27l+1lZUNiZ465ST/93b84K9ipqsL/R1w9ooVKYIKKxCxv5F+j2pf5O7Fv1qhbcu9Zr6xq3nGCF6
Jk3adWXau+E5XyyW67ciV66sybwF/FR1FfvVcQKK7MX8I8/l5IIeDHQiJB6GD3elhAR6WHUL6CDz
uLf6h7cMCSnqs/BeYYQIzBHHsSNqb2M6vOOGrmgEoW5CjuKEGVptU5cw8T5yHrF6Z/hZm5OKO/sL
MsXyG8aF2u7vRxm7BETHuxMKuBlaRc0OqrpG/xx35a/XBh6wTgKBc/EIaUoMr/gv0FYCWjHJQYsL
iUs3rmRwRhEm5iCIIlYtauS/ugVdrEM9s2eaazFAjbqPVcW6lq5hhDUYx7PCO9Wnno1W25JKy/WK
qXLWEkbrwMr/BcRjmYmgTj0bzHb4gzo54CFhaAvitDIKso2dMXxFBmiueVpIZB1LRki7wYPgSeFk
/HTW99vOeHJKrikbv+gl4djIQNBbSkfu/iScVeMJV7dt3SONrIJB2ontlT12qX/3rz286Uq1FSs8
Hab6m/0vn/aS92t296U8Kfz9V9ZGPKZzCHtYWUR0PPvyshAD48WTsUz35u+A7wEnpspT3kbWdxV+
6B0OHxyQBo1jZYeI2RtwAvK/wVtGbWLo8JG8S+THSW9JTCTHu7q/foD9Zaelq70/TDNeDMGv1NzK
UWcnjKd6Zv6Kyxx0ygkjOeNYYncrPFbRkAX5agoK0m6PT/U/GT763XXPYGpU2tGhN2Le6AtK16Dc
86bwJLac+53bBQZrh6qMmy8/t5113RxDuIsxYcAAl2H2AF9ElU5CXqQk8c9uWyQsqjAk3uP0Moc6
T9ggZZw42aTwXp4+Qq9q7Emu4zscWeU1yR3YIu0Sim82/N7SiS3pd9ETqWLck6JwNUvZGvVI/ure
Ew/6qQuAyIG2tYCHShXAANuEQET0xGHbqgLJ0w7xJsTlGemgdXwJZZaLw37urFjXtK7tkSpnaD6g
vxzba4l2pVR9PFHzeSibU0/hApr8m3eiH3EwP/ljBhOK/RYmuAalxkLo9DcinDBkKPtHFKMbdnWU
DBcQj7S/Hq1HroqWoYHAnTXEXY5qAZ7/tgoqNz3X4TQ0+TFQdB7b0H8XIr9f9zGhzH511zq1HP3s
lcE/G9CnRssP+poKKKegX4lZVqWzrF7OKpfSrTleniE+pZ85xGfdTJHeVGtTx5iCR1IuHWz7ust0
Yr4BkOaCOoZTd4pENDpshLoQQim/dgD5hroM6cY1+ZdJ21IzDNR57BJS5HSLYjnmzwXMO5wt4UfL
YiRKTR5v9z+gVHAwga0fVRneWMKkhae8ZMvoqZyTtCCq0wVcK+uuQrqhxDiD5LbuDFbvk/5LhjTx
o+k60d2DPPECukED1UyDg2/8kBUtX6REkev10b4ORvOMVjpia9/iHzumLhXB9WNqI4i4y8c09Vzw
LiwZu00NQ6U5TWYBlO8qo4oZmlZtCBQgIedGREETqTOXEOwQ9xxOKhu4oeFnF755JgMrWx0G0Kpq
LWboz5HwMpZCgrsLMTLkOOks/GBFCxjqM0DlDSifW24PjULh0HXwnQtu4ZVzoJcKo2ZanRODgcuF
XHixdfMSXefpaN7RFDE5gwVxFmBdw0WteUGRT9ke3bnummTSIuzmX5FwYqT7bAGgfjZNimBPT0hA
GSHuL1pzRD0fnvMz6OZ3pqBQ4GADVn687ZA/cbb5lQtUylaPyfXI44vtoC+aKFc827r6JhCcyaZ/
XKOi5jJTanUNEWpVsSP+TxR7U1ko01Y8+k41Z3GYfbPKYqAkUmWKZrZSlVibooPNAPydU7glXBSQ
XDqCYrsI4NLys1dgzfT4pSh+gjLNEnbAV9c0n4nqvP9ejfYr2+WJHKKyBmavbJtYhFVATeg3McfF
WtMXdB44C889OHQdow12eDMjw/VHK/Nz6N+XMzlJ3ySSD+cTyuhd4ZvDWAyuLr1KKK8FVhg+6PXR
TjzYIpjMtGxep7odeStFCBRZZ1yZQQ4JudomVXzm0LULHKAg/k8dgKvLgyiUY5FKBOKHtMh5UQ3V
9FVIHaA1OqoB9rEfyWtgwcmZrIaQf6/QZLhYzCpyzkdgI5CLuqF3Sx1ARnJxLkqVBoDCJEGS+lQT
YOXya9PuANvFm32wZmTmmBixoGSI5NiIL+lllkmZZ9/DJTkaOJEH+x0QMA8haGEFOD0leNCOYk7D
yQW13Zb0H5NJW9lTstiK3Q7N0nTBGs8UeMz3WZCmxEjyDNK6g21lTwPvbXVXPz318OQ/nNnWrp0C
jUpcZdNw8fBV1NK4Vy9rApKa5JHtTSnsTebupq6OddkeJQ8891LGwQv5LaB3Z5sRiPWO6ZBfb6Td
B+VPrvAocnB5YiHmUtjVmszy89P5XphJnfnZRN0I4X49mXQSEN1Dv5Cjc1ZQe4ZZaaulo23XbEoa
NUL4AslWr9Jv2WoAzcr8hd5wwBj6mtFu73AKDja/u2T0pmL4bwVPs5FfO/Xg9OeoI3qpNNRIcDzx
7LkJQiZFB+G6Zqg7oat2Su3QHv/QsemQYieMxgDDnshhCfHQ2N+2rk4CxPJH1+Q322r7xMp/0Zeh
yXYauxOK1pgvH2ygkEdMDBlbIcSAYxOiYGmAHi8i1Fr6pMt+QeVSlXrvUXgMgOj+j2W2fCJl7LP/
/pZe+J16GF4lN5NQhZEEgpcq8NtjSd8CORWzRWJdXzCtzqnMl0HX5XCNof5f5u3iVYgctned2iDL
tiivAt8pGxCgUxk5qIVHspupDNiNP/9R1Yzl1Jveqyr/120P2lEmkzV+5cIa3xCn2pQ9B+aLlSAU
qapTqBzr6CcoKDORNF7yx9IAZbKa2BHRi1ssppBAVvjWXhq8k+mExHASroc7obui0wJLa9REGVhJ
AOZ1eYnNkJIb5qAtVhu5V5n2kCKeuX/fxudlZihE7Xx6WDf9wLZcjbuLrJvHpNnYpFpAWiymCHev
Y4adfFFEnNUoKld6clPjBdaIIkLYTse+SbdvrVBSabGtZ70SAkIDzHU9iYLtNQ6fbpOucOWVVfnR
e3ahLFWAUbgYdsGn3v1RoqcBbNk9QO53SSH80PJ/GgcFkZ77XN6KjjdEGPCoe3FuwmfnRsoq7rca
zn/rq8rvyCRwTDD7osePzWSLP3xYREJ0dd/NisKkQ/uQpA3GdMft5BjJMuqgpIAcSMkO8V3j2xX/
T3tQw47OMQn9wWI+n/Aw+vLVXb9XtW1MaLoP50b5Ch03UzKMYc6c1I7TMgC6qhShSR667R3Fx1Y5
bZoK++Hjq9u9weprptlgMIyCMpvP4ka1iYR3RgkggexMLTiQXJjnl5QUkeC+AHDJlTO1ZT2nhjc2
AEBU6Je/+mzDL1q9y0TD0JFeERb5tAxoLVobxR4T7XCjLmrzs69rzvyrPR/b/B99QUhjpBkq4jt7
2tqNt4pXg4EJFvn6Bslaol6KSU0xBwF3AK/QJW9a37GKnY41j4iVTbu4PIT/tdR6nijsp2ggQnEG
sg4vf78eKIHe/BLgEOp+vRYe88GsXSTrFS27I/0ETkpWgfXIvqaJVFBMZ2oLB+taI9WWJ9gujZrT
hbYnPNVSns6UB2V6CwMiDlcKMx+8ULxxKSjBwUND2iM2ADLiMr807xLpadpYDs+6GjJ+cAUjdQtz
695gl602AWaYqfMQSJ3tXBOWJujTW1kn1NFGA3IYEs4ENgAf52sjdPvpENdpTsPizm4O28nL7oa/
fyoA76l7CZ+xcnH9NIS175UxvkmAeTPuX5vvDbaeV6u2KWpod08luijoEdHf2Ft07qAaTTT9lVD1
3Qww20CKiAs84eZzBByAokGnMXzSoOwMBXUMGFqPCBsFdulz1VsHmn/HVzmSWKNCUdOfgvWC9Ycz
RiC3ez2FxZKeytGCbhXi0136awhPmtkLaG2Z7727kiAfXI9RDNMDllVBZcMXcxwzwo4jlO+zQ+fc
03P77xtspngwoApBy7fkPJKgyLqrtEYeAc8xAuaxt02PdLGsWKJwIe2gTcBLfqK4YbsTKG3Ba/o8
lcP68ygmwLmBEaWT1jbslObF3Vozlao4Nfht+aVdRwBXDQPiGJCONk6RzZ+dFWUqg2svnKfl56aR
NsvPppdJ2mYQsnJbYnQ6t8vIcZLBaAgryaLdjRkJXhamXIailNK8zMX8PIMrFx+OKlaj2n5Ju0Q+
L8PZXQwaE5bJxkcqjjcOzkwU38dZpdO9tJi3C5pCxPAhgjXrIFSkyrLn4vv5Vod+Vj3kAjjRtBqk
iZfdX2jkLOKjlj1D/HmgXbST2x0wax/VRtZisBNi1h+jJXPaHvMfxRRrlEm+urYvhIVrNeyk4p4a
IPkzpLdAsiSC+ayV4OeiRXkC++StDjhmvj5GU/ZTG6OgOmTH8T/pZEyWvPN68uCZxebY7QbF77aR
kRyKAKPPubCaPzKeO5Yh8btvYtjsn/r5bJ/WeveM3jhSjzScUfJWMccZWbG9Qqx6n32NK0CUV54p
X/C8DmV1vNFs4UcmxlbH4PvERXg5emgwEyZ0QrsfgTtGYNgY+oSUwp9OLZdjhh4rT23JIRuMP31j
I1a+M7vPBAu73k7n1f5Tr+BA5K4yFgyCsUl3QSBrjQROlDmD/o4jP/FRsLUmV7knRQSROOIS93We
BAbj8IuHddAFkApx5pmHIjm9NIlda3UmlG06YUtC+3ZX0yerAXCw+i2zsy7agzHEP+x+xh+2aVCF
7SinKiZzur9lIzyXtxP87H0Il7Ml3JQZA8g62bzrq1tD2w053dbz0MnTPMND4niJiXbHmb2BY2js
S0Zr+pvz6tzfhIV6y9muk+WAp6MAujox0+fqlNjjTf1uReAPgP/iVe3XJm6Um3gccAaVzYN7d9tl
kw5Wx/+YKW+oaGyEvz4fx9Kdl3gthXofCjG46ZobQuWeCuTUuS7PxACqKnaSvYhghTl+4+sNsBS7
iLWQ5Db4rja/CuZi6L5r0tSD77SqRl/mRwuIg8mMPwmakfOocBc4V66Bfq9b77i65GKqdZ2yV1RG
QMFN+NFlzVTgn/frazV1QUv3vz4MFXLDz/JOL9fqF4/v1zAENUFCa9tU7tYTFCFKHxaU4BOTYPpn
x8Ba3NiWMCD2cCPTFSISj03zVmg05zWf+0f7w/EoLC3I8jmU3olxxt1KRKLhPJyfeZTMa9F3nFpk
U6ShV7U5OpDaXUw2paNhIsgjnbdU8SZcALxFKZH3phbnf142o+BiAFAr2qg2n6MNUcXjIXcOYZjb
lddYZC0P8/l2mdpScH5IXDZow1NmYy6PkubGtwkQQiJvPLWRLuh/piyLT/Pz6LtorrEGXF0oVMX8
YG/0mNsG+cJf73W+/BfPlqi+dv/ypXUap9gPNn29c36vTnjv08wlEHnTpQR6sv/SFfUPWyOVvWn1
A9CT9+vW81WtsfpdeDvYG5rWygkFMtl6Ajuf9DyTxTj+uYowfZbXQUhR08pM58TjiyyBRZHFuKNj
81dqXoy44HFXkCKGZSCOqw3EESLoA1lp1xL26a9fJdxwJDt/B8jfBmWLcgVUgNq8OPz3OjZRy8Hl
8bILG5IHKgehhEFMT5UIuBOohaLVy7wTXwG2Ftp2pb/vhBgTn6pvNglx9br2w6dkKBt8AQfEBqrJ
v4NODEpeP8pboaX2/WVWrkZvjxGX/8+Yh6NrlE/vHAUWzhM+1OnJz46iy6Xv3sScnuXYXoYszONY
VPHruOVstcwwG7fJHDh254gyeunkAMLOWmSvXNZ+3ne/3yKEWRvm8vEO3upXnIp2W/VauuXhRJ3J
xptVl1NIG1Srm4hyAsqPxFCj965oTVsjp4z8qpDBmqiRSZSQjxhyXuGITo0LbBP6IIT3E97I9QCy
yYTtcPkdgKbGtI/8lIEMoya+NEiqtOK5IMXrdP9JaSBYoXfxITbep0VTJAem6ydmCY6ChBUZwJDl
GByawVzIfEeNR7NbEW+ezprwGe1HvygkLYeBF5TV5avWkUEs+QtmydG/YWAXMfGh3MkcNAQYm4Xr
LDniH5GaRJ6lc7rP1YVgaoKCF57Mrnm7OS+4Ib4nCQh8vSTo8SMW+eH7Tx6UtZQTciqLus3fUNsR
Ta94N5X3rjtd8HRSD/79qA8yP+mxbr1U9Y+MJ87uaHg32AdeBulUyJ2Z8yTVp+gxFOA+gkCEMNSk
Bi7xb5fYTqTqCCC5ssJ++nTzpzHYHGORGMHPD5uwy3DUitONA2lQRZU7jY8qIqbJUAEx4b8AFlla
JwY4KbCX7waLVU38N1X18TtFrd1cCMxK5nbhhsXF+k8RpMMDSh4eMRQQpDQPnqbpS4SizsCYHUcp
n2Ecnjx/5PH2ywdLAbk3clWWxk48A0S4XEXQE+DnV6jW21ZZIBUapy8JZZ7qImfdppZ/nkjur2lo
M8VbhW2uWIGRb2ud0AnQlVHLJnWCVH+KuxJXLQxzj1IA0y7gVFRUX+JpFyKxMH7NuuiIhZRUKpZ7
GbpsYMEuVEEU5cb4PhXobTb3028QlvT+fagSljysyMlNdIb/W8aKYjfNSkenBtO/fheOxvJIHVjY
/JWsuGxFk3bGI9zXqfs7bpsogmGzbILrptv9i76r3xMDa0uBedApoIfvnhGd40KxaMykF87ko61b
cHFk0xokKWft+aaZ/XsS/UFloHZWg6joPXv010jk6tgTLVz4+v7wIsyiGZ/54nN5gXrLnfdflDDn
nYwqgK0DlsowE8tvFTavU6AznFXidgU1IPYXSaPG91T6shyjikIj7QI3In3ipXJCKYU0nKPKFNf4
rjgj0egliH97tTi7hOnlVSlVvkabnv2AUycJx7U4DdBDzLLtZtiq/6+EX1+Lm8diAE1xUYkp8TFd
iF0Q86aOvqhSXMPce2atPUgxj4U/zY4y1/x9qhzqC5zwI5DBfu8RxqqYcGhxLTimLvCYescM67vA
dH3MspJcSTnCK1sOu9afRPLmOy1dpZvxtUlawFr8SPEdorTRE8M03kPoy5rcB5rZYPufB+Na2i1o
oDgH66T19T4S8tB6iHHblkr7p8mKHPC0Q1460htgrvcQSVCDWUCl9vezD2w2FRY65bD+edshEA3I
jTSpvPpY5yT+OnhM57YFBEgNbNBOAK4hTRoe8WVasmjXTVSOxG0bgBodk+9GCMzVKZpMLU3FfA88
CDNYDJaMvOSJg8JiMSHQgh470r4GGHnR82jxiKctuV546BqFYCkqv5J+GpykZQYQCF3bAnR2gxBZ
2WtFgyJxHU/tZK1fZmC6aOdqt5vEWihkd3wCPl0lMMo5W4BNoVDbILNH8FmyJe3pIO5NH7W3HukF
kmNN8HY8qzzQKXUu/4UMcW9eCBU3P20H2qYQ8o7CO1XR3FaAisWNgNDvnOe3a6PPDB6oLC95mlTp
cFQoJK4vXdgwnfd0xsNuv+Lx3eEozvcG8UZGVpvuSIYqrfCSvoeMCim6/HDppWDogt5AiGbdNZd3
WylET+G2mziGm66BDRx8q3Vzte0v4ptUxVYl7bfv8oJFwn6Dt7YHNcu1sOb0JZhGm0GtAXM7157g
LIu/Kj6rz7UMNIIWP1Vdtgg24ZEo+s4cVVcrmfD8cG3X3Wm2KxyCMpUhhLAQZrdu4imMLcwM+dhR
zd49lRTvXrcYWfeyclWRCeNNtXCcjgO4cRIbumbPnsxN/UeKq7E59m0B0cVls1VsU7J7wZDweMG/
U7SEL3WhfH+O9NYAG6a9Uea2/+np+2U0TxnIdGKajHqQkAT2A08HdGmIb5Bz9SXnJey8mNtbILNw
0333sYUplKOirX1ayETEtxufoZ0afCtJysZrEF1X6grL3arXO0OzX5eonFHSVVB1XUW6BPmAlqzr
XEBXm1U3Mn+/VTkEzAIWDjC4Wif1eVESSbzxLa4TIgfymIyNJGUM9noInippp4k9cc/0fMEj31hQ
14trvRVaJqTakUovGmDuCiWoyutIlApSBmh4jsEszswQN0n5KLfJOacF4+CiZawdM4lBpVLR24oP
t8ud4ZbRwePF2O++n+JezX2Jvu3nkPAvgXOF5AizSZxHamj5kJ8FqKy4CyGqAN3LiyWJ/a6U841Q
4q4CpA9Hif4uMpH+yIAdSoa+d+omIZ3d0VL2xq24JuogEJ4YjI5u2dmaqdA0d8EZ6pU5/CJSmKKH
Hwks9Yhz0TLSUctT6gBmnBB16YHG2g+pO7zlYQJQZYOkXTdRTrlt1uLuB5jxBm8yXnpD6Cdj/v+C
/BxRZEDUMspQTiSqD7i9vs1XArvMOws/V+awXBNUVKIvzmsuKWsUJkQ4GpEIQextH/vFN9sbIE6R
ewALfbymfi8m90puydEFU/HZ7oUcDNFQ7xk/bEJOOfbUv0DbmxdbkfrZDT66vrMclQ9bIgta4psB
DLFCc1qGTi4673DDbNZYh1rt8r+wmd9GHx82ma7x1CEfsNnc8QPyJojcfKV7GMohYHE2FF6Eh7gV
Hp7CdTm11EfQrLk8+DE7S6tbETx7xq5Cuc6A76342yYQY5zjCJ+9T3rs1OU5XSNz8fgdahmw7QaZ
+5XmEDUfzAZG9dDMcdnm1QTmBdGvxpWg4dv4WUTXvTRrujKd5/m6JaUkIY/S8/46rTEXoaFoO9S8
AQnrwa6EyAD6BpkjfRexCoPl2nIUY7WJjoa+oYAkSMQx6zHj+5tMd49OGV5FZ0S2rojps7TTl1td
cLflh26Nbs6voYoMlJIZP3SkaJnrQu20rygqgdImGhcBQFCl/GT/V6vFODe8oF7nOKBGKuCGz7hi
WC72k7zK0B3mOOPPKl/tFxQSwwCBvTanfFZipW/XEfjHMRfvbFzNClAo4ngHmSuRkTTVjmDXmTYa
NdFm2qOtDg6yq1BX1RWrwarQVTGTxPDyPZ4ITEDnlGb3ld6FYqNRSCLrF/hXbb6tV7aPYk0ApTFG
FVtARMcAf3+U61gceswCEWSueWGx14gjOCzAIEbdfpvMDTVfW2v4GksdQrOWCIXrTm65w4aEi2Gb
riKn994FRxAVb3rbX5i3CnIz12v/0n2OuPDUn8TVZkidRzPSi8i/NZe3zz4O3tQ3Q7X33DaU0rN7
VHvLyrcwcAl/DDTogDMjySYZV74Reei81sAIqYDa/5LeMbz6AFcTeRpedq0vUirr8d6kPS8q0b1O
9KZnYmSxiybulO6R/i6zTwBKdWB0HHuvml2mweo2+1ei0JomgoaT+OAjvMXlU0MOjTA2owCBwVbX
0svjNDtRwjwImCbSKqzzCEq9wN96lnO8Ne91tqX12j0QxyHowms6G2Ui+zlMGFR8YffpiaNk+h/I
Jcs1K9b2KrtfVVYwho1h+zuyz0BB2U8ZbE2S2QuBcNzkaUXhCmiX7Mp0tpUZCdsqMboM0Qw6t6or
E4iSNM/YIC9mmIR7zsfO7RJFy17R/iwuHF7C1GIWGP4VCKZjXRKrqyUveg5Rhm7wV1uPJmbjdcWl
lCZsN1alxcuXryepEL69XcDUmbmHzKa10d20fL9S4E2pZOVTQIglxBmQD82WUer6N6M2BGfO5T+n
SI5meMuLXIBJX1lgV5CFzDAPRrSBzQql0kouXeNe3uincLOLxU6Xbpmnr+S+KrsQRhobsGfT73rK
ThHFnJE0g/HWk24rxS9gCO6kFqr1DmSivrI7WXc9GS8tR9yeKgUYcW3tFRcxj/l/jSOtSCtabbMj
WWOp9r3zKVhy8u0xIbfcrPVQ9F6yC8m3hVTp6sI+RsK7DtV4JqTPpTRXeOB9xHM80lcOOhnE4BjL
JLz7kF4plHOME+1ERJN2z+7r/eDvEm5m6UdaNickd+mHNrH9RWQvIAnxhuu1rB3nllDmRG3ErNny
TEEnj3EZUVLrzj2yyvDs22sRf8euTf0RNRvhlVRqAZcT0wOxU0f8PIBjjw8VHPq9pmJhQIFfpSGG
MBia9Mq52+G3inqheMDbI+xavR8Ww91dqt0jClfaCLeEjsSWXhOA7UkbwY3R5ff1xkwJ0lUTqy+C
c322Xf+z6brTWiC8TQlsAn5O/yI5GgwjdFN9WDVGZd5XsVtKzGyddfWpMBJO5RCikfoh3y/9x6GY
Z58jxyC6mgJdyLxJ9i1WZdurfpY3CW0S5DOW1uFCzt4VpkcwOHV2exYj1WHEOSoWjJmLLyjGvx1E
6e7vjzIiHxKwgTeA8BuW8uBAEdOKGma2UFfswx1/DORMabxygC+AXh6nOAOr0IkYOzP0WmHBdDrj
HWajS+ZwZO9rLZdyRrRUEG7lRjeY/IYJWrjq9AMNlFIhAR59BZNVxVw8aT1inHCaFw1H0WEXFW6p
oxxCdRbQvFzAczEw/vVFOlU6QUX+Lo2jnaMKEdGnaUCAMkD1EgM0PykZZ897FyYwtIVWWC+O1gtW
UEcyMHRUKUAHOACfY9B5cl1mqt+gJJVpIWzJKi0hhxssd7yuHSJEQyNBdtgVEeaAnHwCFzhnz4Zn
stfYyBItcVxMcDAdrVnv+jc/OGMW66ZC6wIVz4rNOhpQ6+yiwR+LoEBmGKq/Q03AS5z872i4V+sZ
45sh3rcuzwyK7YtvmwvEtltPmgKQyoBkUJ5xP6bGPLShOmKfCe3hyaPIaTw2CMUeWrfGhZeBB1Dy
a4VcyGF7Ki8V4R5WIWvRr/dCkU78Fjt+9CoS5LyNOJC0ozQEDtoU5663sZ1bh6W+ey3ITra+wWD5
8HZ9/9EPNGdwlvQ2iBg5YgESG4dJyQvhbWmCGSDZeDInCZpbAET5zIOZpT6B+PEJuswZ/DnAwIBS
ZlmFSFKqiclbSCCSXGFBDo+dt/AND5zAwMOlPqUVlEFjRhjWBWKv8xcz4FBkaUWbFcgzMJvBwL5r
cUqdZxlG0Q550dd68xNBuqPM/SsISP1jzqZRqmHRXnquSm7MZXVlYAjTPNQwIqJWkfeWOXMX7w5F
kTW9Aq43Zuq3xvjkN8rJ9TlGcKKZF8uGJmopAscK3Gk+XdRsWgoUpi5R0dznlCsOMFdduJzja7pW
lP7vZoOvU+w4tEGdZHfbxttYeOMCgeeMCiPDOfJABKaIP0rN5RALV1gnk4sutLFesOzF/XCT18Jj
oek7pTrF9ZZL6MqpWpeaTmy1hfJEX+mN5SauaUYUUUvy4VwF0o1pzmnGeq6A7LYaJI+mlxZ6g8rA
QAuAwRyPe5G8gvua8/rFCQ6qq8Wb4n++9aS1faC+ci9bDvkQaXFEhnlO2hEJ/GUALWxBMmTugcuL
zsrtcyRB5NIpScViA0rmAGCgMUhpjBWVvg2OfYK0Mcq1lC5gu3E5lFpTqgShLQd1+2E/GyQzpTEh
0QaJTAOxVKfileGtPRDnV1WXkvEPpCZ9MlBMo7H+KGJrHsVpsdJ1/uytg5udtoR/rXRL07vkYtAs
HPH+g8cqtYu/Sg2qe6fn/pnYzAxL3ZL9nnmKWp/3beCzvKx+lODYIXtt9W9IYsKVDq4Ejt8vYUbt
qfDhCnYIjPNRSEfvuWoNS/9M/Nx0QFgUSh+QAc8SeBMX5papsxJBZYKC0HJyfmAOSSqp5XrRrzfp
6mShL+noG+nI8K+Xm/Pf7wKb4i1iazwCQ5wQ45LhuOaaCWS/ic+f3XrecikTEBy9oPUzTjUt+f7W
XWXx7e7O16qJW8yx3XZCFWdRrEzdNrMGv1oKZUFcZoHCkLJGg/xKmawidFvZm/eI24Rsg2G0x+jM
TGQ3SRL0EA7+BoZO8GFk2PE7t+hwaGUPHoPFy/V8CpvaHy2KR5ZeM223t2zYXeHUSEuod5z+vkwb
p8+IBeoN8jK9ujR+Gl8gWmMLgmrfAYnPnC+AAsMGhyqy4M7QmenFJ7iTz9o0m91v70PLiC7WMnyd
jOaUgZINlsBLPknTv3jYMlcS0nk3QEtbfmCxtqpsd7aVSmtboQPuXsvUTeVTird0Vz6E3Y0lcWV5
/qhX1pOa88Cnx191qGi02EeH0/C43wTSy/L48Y14n1MmVKE9+H0KEvtgbuPw/ka+zxl6kZfmhbLQ
iVglrY8iJhnUm6ISn5XT5Sdcj0+Ii4vKP8UwHPXBsOTJw3y7ZXl2SaRPG4dcta9EcMyPNlHihYDM
aoH0bRnJZfz4sCsdYy1lWyauUo1ap/OjPC8ueI4+iYG6+LDOqlNv7CQC8zFXeCTeqHlFgYN0sRzy
edOw6iTpXtvnAal9wknvld27gr1JV0RAFE39/iCwwffashKFSOfBLdBG1HFB+YxtOjUdReHAWX2d
sXVViRN9Og3eUEX0K/i2SSmWrTvv/huVh4cyZ9bKTfA0qtLUxqsbbjzgHHGVlrF246l+4RWCljwC
oiOhnE0PKUDPac7gScmHZnOT+oJhhc2ZpWA9G+rJgmWF+rLxH2VRWlPjR0OAEXEkv005Hg/ReP0s
vWMsogYmSfe4iNW8v9af0e2CaVicCCku4qDXv7B64ydXD8f0jUhBPQkHimH+LSBYhbEV1vOswi9t
v1NwmMq9TqjuGaui9KefGTbggMf/cCXihdbwj4b5PsG3hN0j2f3EZXOIH2bH0C29sHjYnJD3+U+p
qb6ODbI/fEtofUUzJqVr9RgOFdjmVFjOyhDKM2thPeZFZGhFXqI1lPNdI1yFEdKhXWCsERPS6oe6
oB43Wcj572BAOt4RzflwymjRh4Sm9v3XKq5nIIVNQRoGSfWuDuOwMS7NcmechnMa5vRqbpTVAudT
1awySnvXomoc/1U4PfkSY1bYY8tpZ5pB3ly4iXr0Mm1aakn8+o9ZRDs0FS4eVEYoRRwMV1zet2Df
MuezdbVkGEAAFpPd2y/gPOD6h/cXyOx1T1PIp75ZE4jPOy8SBpcVCom1WaPOeL1FclMQZB1PH5j7
32P9M6ith2cvgMfXXq/TVxYikDwM3Lyd5T+cZEE1843FH7mYGS81pm3ZuzhNiNQjAKoqBycJyYtR
3CjBbv8hQ4niHXNHgb69ijP5YeK1vLzYMrFKmskiVLugfpX5pyku0rXiq+OP2b/sfdgoIDIlDVvX
1QpYz4f0ETnzWCTiJF+mslMbPmT0oyK5aBlBmk8vA3ZOihWtiU1OZ+4ipWjjonNqgK6XBCz3HHYg
PoHlgYCL1JGRfDlRnELol8UH/dnX2xaZU1zKhT1y5kWjpRqn2MUNLw5jdOzvIDdC2RaNrCnT6yMI
5tZ8xyFn8ZCqZlvg8fyvScOpENufhmxHTlxefADoP0sUskyuXB+1xe/dFFnapgsVodiKDfKP61ID
pjEp4YxxnfxkQdtwIHMGjSHMXhPslEkuk/jnH76uMtGna0/amQISftkE/SriO+2KnArbR500dNDA
nBSJlXsJ2FyNBC1l07WAmiGUS0zhmoYOuWounDl8oassN66ekOHAi6rggWJ3sv+Sa4pVuntjvAGg
CTcEgVRIMLDFuIM+Ftr191lJ5a6Wsr+nd1bnVTyObOEdXzEs3BfPd6k7dxKfxWn5Is3hEPhV08LQ
RoOAXmIJYjyGcuQHnYZ1JoVKgyITNOPQ9YVKMC3+qL9sBAi0bT3w8ex2up7PHPKio7ORqLF2nfBr
QYKoLUWulVV6NhpQhSxml9FtbnLyFtKhLxrJU06XvC+8gDJj/JrCwt9t+KahFo4fqWY+0MoYBPOm
265KmnqeM+52q9XuhweQ4c9P1lmyqklRWtIBbZTi3TdWofK79zxy6nUgbBLasFcnj0ZmatHmRFwO
svlNao6DMZzq9/nWxD5Ix5fQnNFYBEZrI0PtRlMJxgbW3SU544KR7ecV0iJcFWCtAZKf+SKqDAlP
5I5pE/YeBu6V3NFlTGjVnigy0tuDajGsEOscg0QEh4+DkiITOHio5VE1PfTahY0zx2nWJ77id9Fs
uqidHGXG1LSN7L6zMY/GtueW0LSOgKSuEbLFlmW3F34R3ja9q0vXbfAaZZV9qvZfALDkydVutMRp
zE6Y1FjV+vu5JbKxsq5rXlfMLQb9ZDXhvnFDaoP639H4anUQny/H6qDZePTgbi+1lyFVpDYIyUxR
IU9Jaaop1lG3KLPk8KnaskauwMvU19fFh8gBG+Ojq+afy0k8PdNCWvL84ihgt744hvOgKSyuqoam
6Vy1gAAQekxKRygG7DeCXuUJPeVNAPI0QQ9mKdci8rRLjCg0mjbXT/RIoEnSdd8NqkqfdW492nWj
73uu4DneDjCUycPyAEBYMS7Ayghik0UcNY9druKkCORqh9Iz63rYdB2apbrPE7JtYKb8KdjnUGOu
lbOsscvz8/YTaBa25lVYtJoFJgbLjtnIg3vhhUCcp73JNp8GCzI5fKiAIupVyZ+uO9O5kGs3D10S
f2a9VB11mQtvsJusSNLHix1KGjn7zKYQDd0bHyXYtQ46Sy89UZIU1MgEABcjEkgrhyqaKfhHEga0
JF5GTwnRqqeth18y+KElgySkjEDofUB3mk7Rn3Ll8OHr3o2pvZTFGEkPrm6DmJhC2meNURviqfU2
Ad2Ycky4HJTICNpfoYBR2Miwgy4qaTsd3zsHc/QR+3Y+B9WFwYSbAak1QaOgOaWgyaXTC4snPhzy
PmvQ9L5h7I4qwY3BengBvN9qsIO5dlLBlj6teolASs/CMkRJSHUFBHjmAY5hjZNGAibzWNzMjP0A
EeMWdLqXrV2qc25M4r7925VzwwPzUWXK8FoaK5dCCv2bM4tzHm/jiDtZvs+OwjtpPdLwHuHcuLgD
2bNmNHqCcFfyV6H5MQvO/EVdwq1BvezzWgrNIalfmq1t+haRurevBr4vK8lYOg4uTqO7SENi1/aE
86GSAYMV2YfrCG3UUetD1yxvHJn/UaJ9MI2+rqay+HERfWFstNFdXNBiLmETF9B4Gk2yY1XlzjPj
L/BMgQoOGJyr0cAFafCYWNhkELKtb6lVUyT43ODtS8xHyseI49j/5Sf0pLkbppGOr4xPhpD1AcCR
RCkLGKckjQg/hrhn94Lf5chFpQyi9OQX0RYMSkOzcxOX5Et38o0CeTu5F6cCebaplK2iSmb8xUPh
9wsUYwS19yRmDKGmrNBYPSkagWdTDBFLodJzo1gdF98kW5sCKta0TS2+7wC5ieKavscYXbzwfhvx
b2QDTZWFQycSmjkFwICNfCu0NuvPpyofADf/a1UtF8cmBdw67OwLlakgpuaiQBvXIU7Lch4e0fLh
UPvYlrB9atXvmkFqP4or0auvGZOYZ433GghVhtLGtvgYFLeTTdGrJEhNfHyeDUJfXKdbn27U+P8c
CvZXKMBreCyup/SluD2tr9czDVAKt6iJqSZzzW1ciyl1Pk3LoZdXBBu7DhM6vyW2m2ilLhHhYYlR
ma41NF350IAjhguxiY4zKai4DvcfQwAPdBA1mQaz0+j7OxN44RS1J2ppxH7yNjtNEiRVSXOPD5OZ
xncM6wJBul5wtX9DGQYKkB9FRSg1P78RdtAW4EbYOEEA3+04MAEBq/yW7nXUg6Tav93UWCGBY9Cr
TUD2j52ArHMfgnLuP83rH1PEx2VfGDodNud/Tw7Kgwo3sc0XOdphV9frLnOV1WqGCbgEhbFW5egs
VWFtlP19qiUK0eNH9yzn2hU/EAn18N62SfmZlWWlCz0TvBrvZ+f34diLji0w/OWPbjn9fCcDxcsg
EWoLMDF7WcspcNmwx5U8a4jUsZwbqtBVCE+aJWHvX/pcecKu4zv6f7eyzSXPJM+hQG7rl+/NGmw0
fESavHMMplLGroUmSp/eDKPFrxuxfaEaIbLYpf/PJGSkKGHCox03juYmxXCzQo2lpQrUpWamntO5
fxkBuLn84OmCOPjw9nvyLAf6VYqoiCBjyERD2nTf0AmUWT0HmuhHN1UTPPeKIns/ztUZTCEaphFa
MQhn1fip4omXYnRlj11SoGC2g3/tLN6xM5aY9xL7kTWZajOfmosG4owhaOrJkSfduqLKJu9UzddS
Mzw7ilDTi17JsZ38ok+I05y2SiB16or+k5J8k7nUcB1LJYr7fVeNLhKUmMvHMdLK/frjG8L87MvJ
9nwh2VfBRtDScXVUiIIqqtvEy0SST8FJAjnCDkbSjVT4UlZvq7hpxXZZFCw4A/OHk+su+dzUsFXb
cJ8qRHuxesQ/yyLCbbcMDyStpk8YiZ7QQkHSHv2NNKPOIkpTaHRhofc4F3DzZPxHSKqOUI8TeJ+b
WNpAQJ4x0McdBl65J370J+G0Jr/CUAvn6hmgYUd2uHLIQeWWBPIfwYHFz4DJftuugSaRZr9Rhwzz
bHiSfphGji3n5RUonc9W5/k6b4ZDEGv3+CtvoF/rLMlwB5xUw3k3yl3xCwF91CnzHNb6SecLhfrJ
AHZoC5Vzl5pItGarjk36QRTjH1Yi7nxeSELgnnur/IBHakwgo+0flFyeWiT/g5MBNrFMOrkxZ8dd
L/mzN1rpis1QcMsFQhIEdgU8sgN0HCim+PUZ0lU9EuEWYL7myxyTrbb0qY1EyvLS03L6x/6d8jYz
ciAs8zv/ZYR6/smplIsMBSsh4AWUOrN97cWLEWm0XUMv+uMcNy0CY9UU7vjHRq5p8sC0UBLPRKsU
FA/oEkzbO7cF+CLC7B/sUFhD1tLfFdQl86CIthWdBGko8cMlzcIuQp5uOTLM5OKrCercRi9bDmde
Q3RSWV1TlmhM6R2HMc41tK3PHHgCoOW7b0sRhyLDs2e6mnGfCrKSkOxnGDn18XytqYSVZD8uSh4E
DGVaV6eWjayvEylNFanmOoEQjP2I6giykn8sT8mNEinZIE54dd2RHkuex6ldGiH8J80isLavYROL
VoUyOEMYNrNCioEBMpfDhRJb63FI8t7zmL07jL+/CUIpuyYVyoUI6/zISmfja2V+8vW7ow5oFZS5
9DQJVB6JUvxrHA4jEgnyvVyIFLlCDdjtW3TJWaqsaeoXhmQLBRG9VZSqlT+olnZo6G6JlfFkK24W
ShOOax/Rcqw1U35s+gCWEqC1nz9PHI3SrXN0NWsPvrYMkz68zAfxfNOKL0AUF8StU/73G14FUwce
tuAYZT+O4OtbV+MK4FHYOP4R7fLzRmYKIxPSHddY17+55gOWLJZ2BpI2aIVKK3frETIRSdusZ5iX
vMISLnTDKmVAAcGdzTg7TChO/39vQbERHvWkstJdmOMrxJoRROHh84KrkY94g0NEwdPypGDq2oM5
4wOprMXhU9XRh5IXUsFQfJR3h3NF3YYDuv067cA6rbp6FqBDMnaA9WhZCqV4dZt6ZFqns5VrSdLz
3L4/NGOdYGNtdB46PBJKudLAs6vIhJ0zby+uUFC7J2XUAc+KuHjJ4FPaSoM+bzZHxYGZ+831U4Bs
nzlEVNO2021z0UFtSvJ3I5zk5ZibAgi89bMPxjEx4jyeNiV+0QuTRGlJGLytEYfcnKtrPJVNcxTd
oCj+VOCHUGhXerwd5jEEktiTaMItBO4jzyeudxwlHqgvfW4uGVF+Crt1zVUKACZQDj3/YwuaxFv+
wRf6Ug3EQ7fFLiJ4BAh5stPC2S5/ObRyYssrw9pO9GB3VZUQJi5mnET9fANLQI574oveKSTOLbNn
FZP4ihMLLvzM/euGuPsSrzCvhbM0WlOR4IkPlnyBJ8/G9C0ZJyZRJnv5H5jrfC3k0tdNV0h+nnNi
shl3q5hAXizSwyXtSiK9Mlkd7TfxPGxve0POCmBdxwwTpe5EpKFH5ZHZNuJR81LnfiiAuVFE8WZt
7kXBziZUP/xMURNcePviyYdieV5uvyYmwMUKb3CGm/7P/WxfK+W5fHnCRzn77D79J0M/LLUfmOBV
WlaULXvZ7jpzidw7s8k4nUzxFh6fkUm0uvoE68k1GAs25qGt2vXORB03XXIXXrKCadtVRwLe4FmH
Jlwa12OX0XTMqkaqxzUE/0CVfuma1qPQOsPxI39Zy73c8N83LQD9py8rjUW+6VQG6bsG5wOckHY0
aAvbzohk575tMCg+lTNfEKhRLb2W/o4Luw13ANju/SP5+jSA/Ys1WYU4o9+RiqE8Da7ah6zrjD83
qSXijvvRML/hEQp3Mctwn3Akjt9wTrIUrAAg0hKIAnbuWYJOcnJl2oorCmJY5Q3Nhvvo4rf6YY4j
NOZhuH+vEpty7mQPuVrvrDxzKDLpe4XBd+Qp0AGG4+SI69mFhJP12X7ivqaBw31HZWyqwhGN7zlM
xmgdTTUoXjXFzqVBtI+VwZzguiuyva144klrHVV5wgZqQSUPb7zwWlsLHHhbKxhKKRN2A91YIczs
fsDwDjTgae5a5Vo+CfUXiQD/t1LVJZKKpq1rlVcJyCR8vZyhNOUSwqYyR5nZTkIvsjVFPzFyBCjG
rMK+zNUPLTpgYlYaA68Bb/YB2nMOCvhiMxNZpSSQ5CCmxQ+Q4HOaEvgtMwhDu87SZxLg3P6Nju3V
4v9lWTwt5h7LnuXYoNqv9c4oqtDewXVLwkStPEezRbyskRrIRnpHMbdguMuBqv7sAU+ALjd7xMz4
2tE3U/LKczAEvFI1HKut8BqjD+ojPiA2YOPwb0KQlioMAMFeflROVHWYV6gv3/kYnlldu1Us9VUF
itEgnOif7zkyn3RVc/qnSVNnzN+GkaRsigt/gl0rT4bWZz8v5vxaEEm5m61LCl7DsqPe8b+u+nw7
RFacV5X77HkF7FT+mkEhyqHZFLpoGUMV5uJus3Rq0nxbDZp5CCXgrx9+Fjn0s9pi+XiYuna5KiG0
R4Wt6zJJZknB34HdI39Dz1a7xE15Ag7TmYNl4MvbGidWRtMpeAIbkgOdu8/41v1vFKrKeWiLCpCm
vv3KEcPFtyL/jtd8nwuaQe/iZ2VqKsRKSUvHOHDlkwRPk6JMbVJ/grVvoiOv5A3LmzrPMmEdE3yZ
mnD3I6IY8M6EwMhjppHezv6CUeFypk5ukRSUI1wIRg2FR25+O5S58dl4VZ+KvFu7Gq5+jL9NukQy
BWMNsR/qvX/fRQnahj4nQp+b53CmNU5S5m0RwDsQCTgokDgV9bxKrtChqdkkfTCeUPmOup5Thc2g
CuvQE2TaVSokSX83/TN5+DhHN89zzxMANy3D+dsZqvXy8+BI5Mb2GiDk89MJNk5FsIN1ccT5FdpY
y/US+Op9yNPNgRxIKT8zWTCzJO2trCVJDVuDpFdE8cKLhuhlIAEnkUAX10Sy/sDXaUDp7C+rNJHR
/+h9k/7NFsAmT6lD4Z+hZ5LPWDKo0BF49gFMYxqrwRyebRbSMfp653hRN2bByRjxBbG3MWkkvhPQ
2USKXVVk1XgPa8M/7tmPr8cI11F2vrrPaXYlj40vAu74x8SPXXLXOIFzFGZGMMR3ocXPsUiHXBxX
pPM53IPUX3DorL2rekXLSu1KsLkJx1qPDA/2eeI9Fnq1H/D9wIXwX+wZZUjgM8QoMZxiy0FHB7c9
JldeYbN9u/B7bLUjhHSz5qSEw9+dwujDCRnREB/DSQ49hebw46EcTVJY+eYlJRx3FNsTHHnGtxfZ
562Insv22s/KMIueNBXcT7Eco2ZL5gD/rV6CYUvnJwxezZ5JIvUvPQ/I8cAsvdBRfGESYh82K/7u
9p/0y4Jp0oNjOph16/2Cb5rqRIQ9/m9U8CDXYr9INdEndXdWWIopU3tUyRscLQnREwKXbKj41/Ze
dPmxm/dwJAzdtutrDarN9EMXBKdjOjZJVPLgFU6yQamCBeXXlIZDACw9tZZCB6NLtZVbMezihMa3
FAFkar+Qs3CssIOJirzx0QpNFr77G8JYXnQ3+x5tPQ5qGWVU5iOZv5d40RKVEnuVJUqHfpJBNqwj
eTu8/uaI+oCk1JkDwWztkuoUp9ItuE8bMgbYCtITxyZkvah8WSuQOtzEzcdV2Sp2bd7D426DO1KY
DDi7SnXnTc4SIrMRRiFgidCOuznozWk7yJsrpfkj3gvsxO26AnIZjOr8tPBrNPTJzh9Rj09qatRL
03Ch7u05je4QUzEOz2lmPHsXI1i4wjwRtuaP9xEYj8YURWUuO5QL/lCZta/7OxOtc9tNp9CDF/Zk
engdS1WjhZe7Tkxiq6HB+Qn7lCExp8bHk2p1VZZNTpJOCUtJ3U6i0h2MDPYkBEeMVba1rxQZyWgR
uu0TYoy5x0ajSpGTqY3dljXeLEhzpVGdT8ISY7LrP/6SYfMhRLpuprWU5oMPHgFygaX0Kw9/uG2f
p4BFJN10TOo/YZmwKFDJynAIaKzJLNKFYIZpJDQcxhAkN0OdErFPO5f3smP87YvMWxONGIKC1CxV
C6QkGL7m4ZagBpt5E7gkuw/3sOIbrAzzVe6WR3COrnnznoRV7ukearPqaNomjBQdK4+LYU8viMQS
rU/t3oDIeLSrSCuc+i9QGDvebmbkVqB13oZeWoH//BRusUFR5gZb7lxzJrX63CyS6IY1l2V6NmNw
+oK3UvxzMt0KAEBaj22rF1c3ODIflDA3vzprx96/UsTbLik42i81lqWdg42k622apzUT43QMP2ys
AfQL06ucOI/+TIzji4af4H1SclQNdEWvTM/NClU7qQF4HWaFpDFOaM2t8sjMmsfOUchf3SKleeAY
ToFmWn2D3qRj9Bejg/LNWv9siGSgj4/NAVATVxlHw9Fi76yW1dtnC0W6f7mCkqFhnIIXvAsBMIUI
f2Csv+2Cbo5qDMGpPnXQay571XWS6+Y3ivsI8nazgr68t0+OcGi+r8Gw09KRhYLQihZr2c2qwMMT
1GoPZ4pOE4mQFSVOS+Ab6fnrR8irs0NYt8quKxcTpv80Jr5LovXL8H/4o2vSLDWujmdJhiZAld1d
aT42qdkyYdtkO6QLoGh+TUq4M+p18q4508AgEr20p0mQAv5ou6jOX6wHBi61HKFBeKRyl6vHnMg5
w8SIxgdR/HysbXRWu7495gZmNVBGfPPo0nLMVLfB9O8zCbBIKP0rZucF7afy5gHaUPERxgMHsSx+
gXwqxSpM3Z+8ht9haBZH3KjsS9kBpfnkmmc8InFu5ewioRW9GZrB857cX8tL0y4rvCf578pFhDeD
juOocFUVFUZihjIxCdCMxdo/x7N/XELX+J4kiD5qwbwFF0zazU14Lnbv6W31nPnbFjBM6v7cfFTK
5Jbb+Me24UD/F92JGsz/8Hqqp45eQd1KD5k7IWNqEHQRvcMcKpUgys09OXWB3q4YzC7zlTL8Guv6
iIFLA5G6v3glGSl0tQdiudqf4rYXFcL3/9lJmkCfEzp3Rb0WWixXKD0cDVqVQbyJCK1TbCz3BD0H
QBgZmU1CU5nIf1l8sF6XPCt0zXTepVwvAQAzZwHqGAvVXcK5eNVXM435yhpEP2TBiil4QZk4Bcb/
VUCSFM2Ewd2VDXp4UgZtP97oL9cJbgGvwt1/yuDCKZ7u7LLtwfSHV2HR8hafsvBmlZDpttg+MB4Y
oCd79nTG7BubQnb7UweiiYWAyADJCis6tKe8LnLaZ0rfD0MVdCX+OTBNfB4EWeLGSKgV5uXwpBs6
0mjpSqHddEkhgmI2iaIBvOPGGcxf80GLq+/xGEL/P7Yq547CW2bcM0p8OJg45ScGo0g1DIQFAsic
2ijU9TxO6IkwovzA1r5Q9JgCy2XTXeqW3tVE/SLkNk4JKwKvATsFqzF5QfToaWYA9+7IxGd1GFMB
WTcir802OCxtzQ9K9JM01c+wUg0Ky3It3iZGveHbwNVtONJg7h6npycGR+ar04G3kpfXCc0Laqnw
Zeswwy9RP5Xg0ge0SqPMgXAO/YGY9+TyEE+Z70ERSWn+GhBh8YnLE4cEydHfwbGZJZGmRGGX/vmK
jC2FLWOeJL8zU1CKEc0BQgIkM1a2LGx0US8C8W+lN6MRxA+g+GUjqjtMoBTYmDGklgjioYZSyvm+
kWuKSMI/RB2Ulc94OLLUTCIMpe5N2Io2jyDjlNMS6TqkEyD8CZehmVA42iap7jB5AEw1YxAsIM5W
EVe4O0+SSC6hCpupex6tmDUjY85G1tbxOwm8Jg1qcMNwNEzita6FucUJ7fhWmM3taw4/sY/BB+FW
+8kFpZV/KJgctVD7jA1znUMKHYjbyEFJ/yE0P8XBBDlb+1JZ0cbPRlIBJugRtFccwpaLMjktwJJl
OpAqfKHRfI5rxDh0C6m4GQh5pG0gC0Uy0NULiFbF3N5V9j0uzTVWDBds7tKo6nyNoFQnig5CQHmO
at7er5ZwiZav3S3CcqhCYGpqTWvwJS1TNQdSa0NNufW8S2SfYrc2nHpl4rKCJbjIeXuAW4IfcKhv
Y4xh2OtD0Of4UPZi9d4fmGRFJtbM/5YEtWfIZN+6qXOm4ev0/XQ2wXsDM29Q+QdxNqPmnwBU/IJI
qoua4GNJA7kRGx6eI0H4zZd+6BgHXDtZ5x7hqShY+Pu6/fdEdAuPlVc6f6CAXky5xFIavnoMyBDZ
vI9bZzoMnTeVnkfkeJRmwTdVbG9fGT/6n/SbaactGhwIq7Y2XFbAp7dyJmr3NynCoOijZlLFdI3M
xCmf/2tHEWejs1MMfirKYIU6BhOq1xe1aG/0cQu0YWdirm8oxJj188jFsq8aW0jpdAdUfSrtOnb4
jPcTk7uM12ULjvXXKQkfbg17aiscwyd9oAKeyBOT9O3JzN4ZOzZO0Cz6+5GNM/4aHMBh4AATpuif
lRyD1ch4va5nVNtthg6asj30oDhwVCyzdSfxN+dNcQq5kEOqcCDZzUk3hV6OKKliN6zYHAm6b5ES
OcUE3I6/NvlHkgCTP7uiuud2xp3hmjAIuD1zElTM1+ms1EA1TSptpt5RzoFe2oOADuggxyYSBg2e
s0XGxb8nOhrbs4t5tx52Z3fTk2F3aJRk9gZWODSTJ+tBvcIad55QBGeBjrSZB4nLoXJqzDheus/X
CHem/RnO3KGHn8lpIAWQYhBL2bdd66ZhExiwHGRzGsQFPDmOX2IIe+3b6WNu3BiW7QkULjdSDcm3
Qv1j4GYSMZQzO3/ddL4DzmrDYrMG9J7waIXcBM9PIZ9WMwv1KkOdgR2RsoiD3h0WPv1YS6RIwli6
MMgIPkP9puvXbQWrOeh4qGVRX/R6/MekoZLQM4lXALDuufrOIqbagos/ovcatl8oHYJR/DDozhZb
JmHtEmd8/r2xaV56g7kh/U2DEDJfcujcs/bBhs/oDjaDRngyAYTMrk65cZADI4IK1nxoL0Sj5NCe
JSqGuk1SkVwERCXfuYqMyFw7nw2TBCsmwYOuhhQpiKV/zgwKKpBb18IjnE5b3EtLCMD9yn3HbRgm
Rt+FHGmR/CnTJ6vPf13fHzEupzNvo/dUqzeNDYBQqZC49gzGtbHYqNeu8H99teRAY77iF68ZI2wI
l/E7lPddlpTzGAmZu/ZpuYXeKxbcjINU0mcc9zLUFvDJSBZgPX1DCt87CoSp/lqh335SPLZiF0Lb
HqJQJy5047DWoTnF3GDyN6h2HoL28JI52acR68daPEjNOFXyCuVuqvVDIdW6duM/HQNnaSKTn5cY
U1WvXj+BheTx/+U+mkGZOKjwS+JcatmEyp1EJHK4Q55GQB7ihSW3Yx6+MzewZKQY2MIsHs9wdO5e
RtS9ymX95CJPQwVvxY7wN+l/Nc0MBv5I1iyPUcaVYFqML98n7zycXvBiUuBBE1oEtgRJPpUaVnnt
vEHn3NPSAiJ2532mwjXjmt+YZ9SBjPOWwY9ERHI1qUfyVnEnS6U/2vEVSLSxeCLamrPC2+jq3wNI
5V5efcCeEHDyDYI782pgoYytY2hr1+SqGXBUzF0EBWGbwaGscrCywJ1PUa7TVcq1e6gDCNV73qOn
bFBW6wclQ2xR1WZKmYB4nosD1xf+C+vQGE7ydlNloBO97DpAtr10nVEKvpABJEBZ4ozm7PGXeAeJ
zwj1+UC7XjsrGvauGcUcnXhwBZX4ZfOYV9X6RV5tjUV5LnZLKaLxfR1giJKDTkAfMxrAvelkIWfB
+oEn5U1fZGPVQkVYDHkcbQxyYJ8zEBecyLw/YGSmImYciD/SvBPbTnL0DLuaBqADQ9OjZ7Qjl5SB
O9GyPW7ptQRPHp8s/KC2zvEwyI8qcYj9a5lPUYVfQ28ruWZ53Y/Yy6lB6BwPvv0vLz+4/jzoZqEN
Q/yq9/SLA7ZHhXcXjam+/RMb0u4TX44TEGRZ5v0MKzdUbG2E1OuySrZjiCwPRq653JpbYbHCp4Zy
UTxQOGE5aMes4KR4Uj6FgkL9kjStsKGC6P0JnUWG8VIdmfEnx1toBfw2hxLrhd/wH8O1tSLXPOeL
2W64bzZJbExMaYRP/0sPPSN5sPO+6+hTWOiqQHIXqzonppdxZAe2RM0HG/VNV9slwTyNm3tc96hw
Tjkycyjq4zpMy7c/BvzyEe4uvmKgTbs5j/SLIzj0lGPY0n3uCG2C/pvSVLUnTZVl7JRKyXgBmlvy
Quhngt2SaCPrjValC2ray5xqXbR2e9BleqmAJnYYN6anrccSpazqsspSEJYh7lVTfV2ybpczU3fM
5R2CU/HYT87xgHAmUZc/5DCuPCLnmoqNEYoVr4QeVbL/oZp1xy+iRUVZm/9aGxJZGfEs3z6Btf3B
X6GYkebyhc26Gy7H2kqvFO2lCNaBW71O2CKIKdzhp1BS6okb2/x2YwQjnoX1hVm8wIdwPOdSQjKA
YH3MHG+w5b5A0lMsR/IhGxG4FgNU7fV+poI1JvI0TuJCgJ6YZukpH2EKLdN2SA+eYkaLfl2lA3eC
tJRV+REUAMJmYgf+zKvNfGZXjM74O3lh36l0T9mc635p0kjBdcSzMtTRxuruezj/WKqEKJPVX0Io
LLKIKgsOI3H6dOV0qIMZpKNZjyoq9XOYfK26OCkcvo1WToy0rBoUwrI0RnQGy4W5guRdmjlx1Fvg
gw8zk4brzNItWvclGMoqm4v62u5PiB1Gh24rGBpkRqFEvw9L7lAEVVumdJBJIQ+8/51FTUtX+qzV
h4RIcjvFaSOx6o+xWTFmhWIUpKeRnWtpAOSd7dhadnrcMBtnK1dfExOg2RLMs2doBPo6XS/bJcTb
/W2DIYrXUh1246CQTFx0adNPhu7JqXwIv9vMZe79rl5utvxVsM1gphyqQGXnj3NjlGisBcXia/qw
l/hQnjT0QV/HyeQ+E/Um/fQgUEtLZJoafXon7BhG0mV8uyKYhR+uOboZJKKm8rEMFAuJiDNTDRd1
zVIUUF71T0i2W1W4R5wDGx6VLDp2hj9A2DdwriemefQvOZPq8uyADYDtABcscJY1KJDFmAOXLmPB
mXLpyZ7Y7wARVgRT3LdykIQH/NQgsYPM2loCMukx+VjKjwsF6vnUPD8PnFfUD2RVJAbwPlJrNQ2s
E2tIt2fpy0ES355rLxWEPowWso/ky/Mm8WZdHLuC2Gm6TLekUTrE3fITrjuSwNRQixCnp7q2zOvI
wLwsllXZx5kMwtDxvwrE8c4pjfCK/2egzM7ifwSsLVZENkMm3EsWx3JXJikmme7XNR5lTh7ZBob/
UJK4NCqaUFcdyhgrQ92U4ZTATWvsjAf9lNvTXb+6Vv+wVapRffQQQhBdFC0e9UL6DBch6JgffDwa
nW/rsvN0fI4a4jcJvIKWjyrwr0/Td0Q0ut3EqRZtwbL9MFVospN5jRe8aKYTVXR3EnrJh9o7/fHb
zIV+NCKlVPJgpaI9qic1wLo6P5lrDfeJ+JshMG5vYu+qbMpooi74o9EIH4GbPPjkaw2bEYy9Nx8X
iU+dqgOIDX71kY3zq53egS1GyH24Sp4Y7r2grNhZqnr5nP+o0Qnsn6OD2ryu++T0Bcaf8ZzslnG3
qD7d1CT+xcGaFHSXOFAoHLHU3iy8HHziTBWUkjg0A/ICK9mzZKhY/F1rKbn91uEXf3AtbK3GLtmH
AFwUrdVqzgp6rhG12SDwwrUfcGFROBMLZS7zGxDfraOtTPEESBaMzrxdmnKHaDqz7/gvSBdc7N7S
wqLlu86quABi3URHE6HdJQn3DcZt6NKS4jCB2RZFLQY9I0mk8NGOcHl/8RVLMKwathQGQrwfO7NV
qYOFD1+81sDiF9zpEzf01W+GldTGYBgi/4DWIkT8120vJ/11sLsoG2bH1euJ3NfUY4mfss3IZDAH
LL2QsQjKSXnAi2xm0Yd+i9h4nKdyaVYvhhMlUFsq21jbFUZ0zPh6iyhtq23NL11U0F9HCLwKBnRh
iBrjYCeVQ5pYmQNCcWnmXHvXu7WH76y1RrOB7uBDirrJEpjY6rIcSwdwphUlTJqaO0Ri97deK0Sh
FSlsmY6CUay6jLUVHpYwmKp331C4zazQpt4o5q0WZrZCNX7dYoPwll/V2ZogjcNSHCb3JGZpE9Ku
R/LkAXg7fKI1O2Et0BM+kFLVBlOPgMBcUfamILXtSPruVr+XssdHuD7jKV8Mqw3HR8fFEUN9n5NY
rglwIhn0fMKiLNwKja//TYVzCch3XIk7icNEDutAwKNLkdSs4MZyyw4yu3AVzfI2RinpSo5FP8E1
vSx0nPuLv4pUm0Z9rolEPHQ7Ch5PR9+fR/aheVlwtRbvV+2rhhobM0h7H3EtGeBkdxstperd25Ts
B9GyyRKb2rHDnsIq9LP0iNAu/DwSgEobHnK5MzS+0DcYa9Mh+RrkSxwChzMFfZKrh05DEh54/tc+
YwkIAze8vZrczaDHWJE3vWFv483ReTSsKlcL+ZBfBrIo32f489KIpKn1glFigzUQc35DGBEP5RTx
8zyif6Wwb3FXelgON9X4um14356ICTIG/dWvDUjjiRABCjV7nrkYgByUQgao/uB6gH4TarJ5E9fI
przIlFnVKld6l12KCV/C+/RHZJQGfoNR7RQ9DtemAhQOp3vL3AamKdSGnXOigpfi/HMa/CsyfEji
QZ6C9C6tukwftSmPAmGRHg1humu/qFLHhM4Z+104ijmqvVJXc33jHYeoNiLNechLep9uKlMApkDJ
m9MgC4G6EjJQGsXdXepCQ8fUN2LamDD/vfyPhvJ5P9YUyxaV45kMGdPUIkJgkLudmBCIl3mLo+65
JPj9SXcC4su4Q/B2D35RtfGipTdbrMzcdxuqdaRftC7uNwffSvrwc6AEMiG4MS1zg41bs+ZX2gCB
E2DqP0wIXVM3X42t5dOrYwVzWleMRv2boElSQzkqgOLV6oMaW0yeOA+haAAW3v0wm7G5VLxqppuL
fjuSKx26tkaxAxbaOzlG1A61gQdOBsMJSclpzZ7gW0lKNm372TH4kINy5kzUwHgwKFGhWz78WURc
h/DosXQHdaxy3cAIeePTnAYd2uMWF6h8XmOxttTVDAmMmT13q5EYXwYN7PFmm7QiFURTwk+0wHLc
ggmVCDXK/Fc5XaqrSdpe1OAPDlWab+L+L+yXItu7apmGFVYJHsM04SNxbfmDfwWTRJ3cMGsP5m3y
xlvI/i12NgJlld86yScXjqtKsGkXiluR4ilfhp8Bxukyn5sg+daRWDjF9snoKzalPyDfZIkunFbj
rYJu0kAygYohhrpuUHi5rAOmLyVM5xeKYXJ7OPofXB9KAhAdPdXkVGErLWkIB2lrepuIZbPJqdU2
QEPY01cjgo6GREFLjVxKpT4k5IESaxyzROJ3NWuaGmxuiSyDQ5SWkdv8JwwU+7oN5YnrzbICQiUF
1qdRMexhh8y+K9HlrN0APmi/bYCXsJKTvR7XsKSaPnnb5YZigss6nTFcqgvojK18FypA46/6U96r
nVgQXQcPlAePg4B/yt5lVdo/jbB/SJNWxBCq7BNXu6sT3VccTvWdqushpdFqqe5DXUrQ+G2Ai/PA
KQ4rvCIIDs7ReV8WXVZAc4PLy2MSD71B9/pmmEScXRKzUBkPmRwLFykFhmiNfupNw3dvdsU/Dn+0
4ZF1lnQt5krUXpBnhR5Y8fYgktLuOBYjnYOqnAr8ZpQONJtUFg5O9sU6EnhUkTOo/5lgkjwOJcWT
Zx407TgzHVdWdbmpOaBmgM8/BFYI3iQDBN1qYweYLyAgxb/pd9Z0MxVv+q0rY+md8XaUio38gWsI
EgRh60TdSPBfdU/bTnSxWaPYU4F5sH83OPCpJBp5E3lGlM8tc7QCboHXAHrfWUbAonFgRF2Cus82
6H25zHx6spxDUXXWi5hOi7cqw8RRyDOcMGnP0OnXEzrNpI0GjrNLLE/blU35VB89qj6x0NyKbt9N
+3VVsDIBbghltVZo2MjueKFKQdcb1LEmg6zcsJyCiHA2LYyLYyD6RxyXx7R63PGhic0Ensj1Vi6p
KjtuIAUeo6V8EACzvVzyo1OvqJ6LOsubAvY/q2ejYjXdQQ9qMrZJ57hBpHXjFfHAZRsrvA/MK2ix
1Vim+dCw05yj0k2EE3286rGx/BcFjVqYsY+vrUFR+dEL+uIZJ2+CVtkevO7lV+obnGg34w1BsPBw
Zrwwb+JYiXqhpmjvMc7QOsaEdJoRWjrMGef925YklUeSqFOYZrIZiUHkbNT1LSgyRcDcYx3QdZnO
DqKrzP8Gq3hHRPGzcQ6XNjUrwtNPxy1khsxtD8bM1vLNeINpXYtJAucJPYDHG6ch+EtOOpIRTWBO
C+8jap3FNaPwQJZNZvL/eorWcD0t3KUZuxOdO5YWHDAsmH8o4R+Rcew6RZhBV7+nHnsO8KlMTMjt
AFMmmwNO88vEBbRt6X8IQ/iPmrdy4K8ZalmKi0uzjMw8vK9F20z/ZpW5XmqGVn6mRI3F2tKToYJJ
aVLDt5QCqZu88txGfAy7OjcOhG8K7KNRNhx/HycXbtP4xsKPWD3BLPcLZZAowBbqilctWg9oUA1O
hT9J9NOH7l3dAUprN9r+t7RVkhWaTJeB0pD+BixklgS6RsYjS7+JMondDYuLcq2o4mRzTpH479jj
oGEEsaY4aF1reQpCDNzC+qbQs15ocF9nDzNegirMr+IXory2RgqF8cKqNaxu4f9r51t9uggK5YEu
u8LeSM5aVlO8xeECxmAGZNJV1hRSek5tDY7du6ZfXv1myqaD8PVN9Nkhb9+YTBQyFvaoLIYdZavV
ZJxd+Fi3JzrU14N73fJ2VTGT0teCluCRVx/vGeevC2D8oQpZyGjoz7By4k0jp3MrDnh3xJtumPiJ
iTA0+I/m9Eruo9osvGpa+SnxGoVqjsW5rA9MU9AqdTPwQ4CMreBWImsa0mbAgkZaLOvfIprvb3Le
7XtfrEMQwD9DhEyz21aUs7vQ4S4uVhNj3Yucs/5UV/aKLX9FlUZz6vUdvc7ynhQioHnf9teCmfoa
eo8hO5WsC8SjkdB78wCwQAwtRHrKgvEwN7CpanPVyFjOvvFKx0A1WadcqymmuUqA5kmeDIwF4ocU
cj5BPW1Q7Vpd2DlzFGA52dKIAKDSqASGhKgY7pWwMyDUrzFeMrfGfVoRupR5y7DmnQoYB5uuWB3y
Yuf/6na3Q8kJX1S0P/reXRJs6XHF4uDtaNxaprdCqPONZMf8H3K1T7HTOcX1FZDFzmOO6GycwQgw
PsxYUWTmBQmsJndYcS419fs9Mkwp4q0LSy3DqzqICSQjR99Z6AtLXUWzZifoZmY6HjSdbJkgtJ0x
ZRPOWrJIhya5obTkfEbaHwm19nEeIWt7J0XufyxdQB7sbZJnfVziIhh06wIObil9UHML1Ng1DmN8
0kbb1lSKhg+//9xVBvEfynVZo1uDiU6p43Kf7kdcR8P8Y7ZzLmIsQkQ0YNJD6iwMmt4s5Ys97CZj
jatn6XmTgZEgrOO23f/pcwzXCGqczwjhW9PE1M+DjiZyadpKoaQpHukvFfOlYzKseRSRyfsys2WK
8uvkDQHn3bB5JXWXbCsA8CBH+H5UF6mFC6/6LQDqlgWOTia/ocN2VgJy+6MARLAlsQDgAQJ4En4b
lJFxqbC9rAJ+RHW2anZDDNOM4rzrYKkI5kdBsVCWjHaq0V1Iq8m7n+GwSNeNWklFTsQRsa5oD8ck
QVQXwVawDE/C6Dw40rizkARXb8d8pcGQ3xV7IwBAQBFb+nRn/iOEnD5RL+5U6j7T+qCsXfK+Q22F
aTbVwOziiPafybiThNRE1cNJR/+nWPkVnDQpmwdostbuKRllg/fWr4neb0CLQEafqbijAkVxA0S+
9+YzZ2P0BO0aYt0ZiybKgg7v/cJgCRog60yhMGSm6dUjIIDzE98sn5UCm3S7xex6pguXlZQ0szN1
tOuGdHGl2f8Rhsr+LDKt/dW5JvqPF5x3x3YAqCI266Qej6ZzZBaToWCbkY3wSoliwc36K4JgL0OO
fHnh0oGElBwo8r+hUnjcKnBtk2PingVF6ofIudEpc+OkCJYpLUB6jROUeJSYtzZeZWIVOD7qNt2d
y1rzXk9CDR/ZdaROwQlW4491TP07ZSb7EwhP4Ge8FGYgwA4+L6eILU1Z4EYdSEj2XktOMCrGIFDW
R8d/C0Tay6UZez5ppPKQlbuNwf6WpfZEZZv3l5SoJTmyKa9hurqTh1M9qq0sKWKOp+mcHVHle/di
EiPna8n2cSmdLYdiAMe/iQVtL9g7YfFTbdMRvThUy+xm2ZL0IGNjzI7GI2EEuC5HRSXjS57P9Z/a
RpprYU2JUdg3ayvkgPlp5ZgpnkoNs0odGaJNw9FmfQI6sx8HzdtvcGI+6Ugs+HqhYWiivtweU4ov
jqT0LZ3fiYPxg5gzNJC6hhCcPxVoOS64Ckm2lWKU0boR4FCbrlyZw3HPEYKVEDp/GQeudJWhI1bc
H6kJ4neBMLGe4Kqojwf9ttQYe4o+8LKvS1yk8GGEMa3P3p5ebUbDii3QEyBXz+ym+9RL3N9CrmiI
IBndP95XSTtWqE7kqj8Qd5sYuUpLkachcbX9d9VNTp4rUdyHkZ/YbFzGhImuWgKI/yQEp+m0ebph
b8aiKFTAbE/ZY8RkOcc1mn/3b+RWM1qGsE0YJtE0jKWd09DMbxjEQGgD/QIAxmFN9PsURmvpOZeY
5uwDfA8KRT9x7bmaQbcT2NGH0HUVxxzNVKW9D/4au0dAUXx/3YQA0SaSYOSbI8+HlugR0SNC/FXp
8swZusyZP4XABbfcwnLw0ett1hgVZfkcoAGvwel21DmLznarKaf+cf1eB9/eZPqKzDhVCRfMwre0
q915irMUcq3TZv5oreTXfsINZdk9TSzndB3ETsB9N3xMcOOZa4Uq/TmKAR9kQPvXvK3EZkeDjXWW
OEBsZE9vO0yWuqUL+8Ya7jo3fj0p3rHk7+JWpsU9UonBnPzhMCIWj9J5P0vbb9PfsfvUZBtJg74f
KVdaLQx2NsJT09bamn0MGbA+qbn90ASzbOCHhy4pBPR5QS2aDxpV6e6ySrkx14fyaTdpZ+zC+NWW
r1HEgec3mUzEecjCVAqjAW/lQhJfTFjSaIaQRtPVKtiiLCjBNSSXfGMmLin55uY1b666qB8YDfA2
2NmKbkGgC26RWSH4lPr1CkImeNqjMyGALyeXNot2RIyeVzXfFtXll331Vd1H+7RZWru5ytyjDY7j
m84QYesNkpCSpO629UfJwMTAhSkL7FmUrKLWnTxqDMCSBToLe2VxRjp+5v89drEVurWKcpjjpCqv
YeSf9QEFoGj5rZBCGXDH8tTw7cfb9MDFZEWfH+ZIvd8dqM7v+rHAqRQmpNMcfxYsGIHl5/0yC5ja
GopZaYd+Z2s/WakG2aX1Gm7cnkJSupw/HT3unIWscYNm4Kno69L0VcS9TVNLrA4YnbdGOzsq1KVG
GAIe86d9MCKumY8lDY0lO3TmuxH6qss/y2JOFzgcbN6uGYcAiL4sTDJuoX2gGFsUSYMB0TPI0p3+
m2WGSb44e8UpvfMvXawn3s8SOXZdFz8qZ+M5vfP1dtXLCCE1tcEpFWOpVIcR33YtCywgg8IrmPhE
LEJLITEqh2KsMOUup7Vf3YYNrzOx2zk3PP0Z1U9TFAwykpP9NFJ9tBlXj923ww3EE23r2t1+5sM3
doptmQOraRMKgPDVZ0f+hvjCPBnyXTb8Rfoc3KYgPtuo07lVnVSl2rZgpYskq0WqwguQps4h5vmP
BcJFBRbKFN/1htABEEUGqkaOE96n363tqiJrB5owrlqI2jwfqVJmFSWhYAt9/iB/8JtBJH/O56NU
nTH29VwRbUv2zihS6EHboVa1r3q8CskBoWc1MMGVsq0cT5fPKYb65FNSW01MY2X9RkxotXs81Wp9
66eVsPQe7e9eqfXppxw4pFnW22bjHXpuiLjfv+836ylYqaCHcfefvOdyoLfIn5fkT0cnIpeqSE51
mXWyElgvRI65IupogRWdDsW6hLNsPvB1D8WkvKzHoaq3mQsENrze8oQvi+x63Q+lv6VByB/9/0/m
dOJSNRr/lfsv8L1Ha5gJQBocR3IGVH94W0WTOGLI5i6zbUPNKNbubxLeBGefPkc411d0uz06Lhv/
ekDPzXjxpgDO9dUFJy7iwd/qWKtpQ63G/Lb1pzC9H1nllvq4cHoPC+GVSXDyl4BL6xfzV6bruCBz
MrnrFxSBlWWP16Brkl2v+YxUtT2ERjDJnMNyMMprJXe8EsMRpTWwhPXnbhlJfEDFT38f+79WfKdn
516xK3q+N9EK/ZGgI0QS39Pth/kb8dJQ9usPKi2biNtreZyAHFIDwe3i672jU5wsb8Pe6tgnkYYD
tIaG4UZ3mqe8vmfQn59MY5FyFA3KRrBh6N2K5cV4l5bG/LPPT37pwjZf/Sc86NFluzxxtDWmAXKV
kd2Cqx1dBq2ijqoSClKcOpzFx/qpCacWaF5VHLD/vJQDAxG2CXqB6BulDBMIqAAJErIq1TowliGP
/N4HKlVVpmHLGlNdQRPpcblsvrdq2XCH9oj2YLG3L50RBWpagWtFGqo7U2iFQg/9jCW8Ku6dhDw8
XD5l7In6ftet59fwBuJ1UIhlAhFFkPGysoL/rErWtq4ge2pVNaGLlGxIFhkqLqTG0PG4+pzR6/kM
AxRvTqONrZ+mMtpNq7oy+8PmZ4YEcsdqMfAeYSpQ72pbwnRGfq+OBFiRl+3jEEm80+b3R2WITl+a
IBe6HjUhkKwJ1TiDiQOb52EKsr3HsDB8gUINACZcOSm7JevFPaQZu4DJ/bJhWj36ZafDnsMgoOsu
GvgyXiiT5OwkVGS2RIIsI7bLpiB7NjIH9TdZvvLZBb+lJyE22QRUdCoRNqVOKjWI+AFuOvBHuRgJ
CKGXJILrHnZnWKfPcrPqNYVZtgCs3kKgmHO6azMcJkztjwMp0FqLPxjieighnnbEyOL/4VChMzU9
PTSsZSdYpJlXiGl7Yg/eZfxR/C4693AzY36gIsNfJvoIF+nNFlMZdbkl36hKDqG3RjYLaoV+X6er
mCR1muZ5euRptwcaKSnb7ARau9b1KD42o2hR0urWlT81O3B8vyOZy1WzD6pLnIDtECKh5H/ptywR
hZZe+O+86tk8sSbBLvz6mv17IPcVDKwfPlXHbY114d/V8yzfbshXf/pVcUVSjFhOSRytUDgy1BGS
3BcvQzwtOqkcFDXliWyDGkCtNDGZqV7TjEKgt8cKP9oPZ4wduo5vCWKlB2SsRTDK1Hvay1MBUVl8
R5jzhOY/WIRYLtNcKqGlbgqvA/Zx6oh79UFxgVc0NmYe7a1PWxWtneArGK525lWGtygiHLofe0La
v+iukI4z9RMxDV/56e6l9rd7e2jD+cdJPDk7ZSaJhgLHkT6Dw22fQSslj3n73SXTpJ1TO2pZcz0y
1gfat2rJoFiPUHqjnlfcXJM5qJgXcji0QM57aZS4+6fcWYVkpacuCbTEvPom0jROPtuEdVqKyayP
q4qrN3vZRaM4zSJaXAbyRMbuJbSVhr9PMlmm3YJ/6N2LychYQa+hrvqv3b9euhSdjSl/Mo4xrQFj
5bKH3oZhaTFWObtPA2GSijsInCPj9owed6Nw1+EuBBuZkJuOSd3r1RIvOp+xZ4WRhfwt4YvvZNDv
Rz388E2rLzZKTCDoxbIqCrcYx08EvkeWufuWuv7SzvWi74H5YSzKJRC6vOSkgbWAk9NTJ9BIzFba
MX8Yr3nVzvniUbNxKqvw3Ojszb3jF7GneNMg9VWDnVszW68G05fkaIfYmSzpfUYpE4vBJoaadfcE
2g2VrPugbbGkMI+K3Jb9q85Y3TmjDevQy4rzXSJhGhQBxAMo8iThaoQaxlC2UZer2Ikj+Cuj77SS
PmsBLJ0z2rznR6gq2JN86rtB2caZUCGLMc9gkHUi96/az4ALUElXTUkZ+jzwvuBUbDyJRZLXZbUr
tyvabQrLwuVDTHZIaDpUgNdAp0tfMTkCJxDLFpVG5Ry4VCwCTlHy1kJ1BtZ24VdUiehHxQJB5Xkg
+ZIrJ1L0guVVORoza4MPC42D/wZnX276O6SFpGnRyPajdjBVZqxbqUeOCiDERsWBr4UP7dWooeto
g8Vo+Alv/SOe0mSMEFs9/h98tZ0Ukgphp9CdiE7iX95OoG19G2erVMOES2Sf4PwH2/bvYE3nu7Dc
MglbOB5v0pjjStkjhxUuXcdrPk9BMWx6PVx+7KsOLwhn6Z3HeGdB9tTaFEb1fY5I8rnDv9tvSsIK
oKhwdKs13W54AYXu29KqoOrv4wVZ+z7KVeUaGAKOfF0lESVFixNeVoopB/isH0FbUA2VfNX293Z7
YwKVPppKZmNQK7PGU+tSNK9dsJX2LGb4tyV7nJlQ6WPDH5ZrV1tv8QsjxNJQn2wckkm73qXLd+2g
z38O21jxCJvCq1tai7K1bWmLOORLFu5weE8we2zmDjdn6575zj5h7wXFkiXai1fGC6ta4npaZMQk
XTkindRlIuwsePp48Wal8y6SEkIU9Gj2dznVnf2YIeVZB+ga7H8Grbhci8Y2wwTfONhC2m1vJ48f
yuNP4tJtRpAYasdQ6zeqz4bxU7cw+FASYszZ32fkLtFkKVAvmd3mBNiGqe2+P4BFlxMtdeF41DcD
lANgn7I2uznvOkIam17hyV9uTBGH13P3UbXHrD27YsOn3PBEFW0GWXDA8gvwOglVvySylwr+GF8e
ZGDN8h1qOEp50MkYUQOV/wRT/KNGKKZKhpioW/QWOX12cbVcS9abWMwQzszeao/yOK4r6syFwHKf
q9m2wMDOy8rjDfiGQzliPHvrsVakrKGt22PWe5w77LdghJtA64jFjOCLQmk2H0wlQxESULqatJl8
uTMMB67NsfeiB0uvxF84g2aS0xaPCsJwBfNVAVgrSnFuTvsoQPutcDawasTwipTiPPDIMB2a+IfH
wYKYZRPeoWWtBXWHED1QE0fSzd3mLRlcLMI54FAJXIN96c18ZrtFGZJ/u+NC9FnBAgdlvPBLmnf1
b6QhgQ2qtGsemijifw/ct5MMQOInCBaFXlZrsiW/REBZbph8qhaZFIyqKCtILbl4h5BiMmgS/YLm
bDdN2xcdfMIrWI8n4BYPRWeX0+pXkEaVb5XYrfp0o3CiUUx42n8qWpYCDqQgssofwjbd53sFXKj7
ZtmyFopA5JurUMExpEl46DYidcO1KlBFkeiTveHYFHDnR5F6+hEZyALcKsNSsCTlcw1QUtFiXncI
ZRocXK3wx36L3RFXmzi11wmu+n2Gqvd4qzR2Vv7nd8yRRZRsIwd0nbYjaFVoAHCBXfN6lpJ5AZwO
byZtndSrGpi5s9+VhM2doXZ3xbX8CA7VG4S8Spkt8VULSlD1ELF/koNouKyxpx2wtfI6mXaKJFlG
xEJsY4eRuGjYQB0Owq3jh6h7gLIfyyT8MqjAhWfpuvy0GGs96jwg1V29WN3AS2pT02MI8NfeqU5h
5ayEbuyjQPOu6+b7Eip4f6JHqhQNP96hKDveYo3piGRStUsyLff/vgL+xNuvLWsw6zomZVeFgbfO
AwByPiDS99r4M9k6ilFv0UQPZmCdy6rVNEt1hVNHOewdZxS+L5aICxHfoJ7L2UMFQDRPWJGdN0b9
TA2vgNd4ozgv7jNZSOHFKcK9+UZvxQ/MnznWpKLYP6y+MAbQ0kjdQ9K/feIL3Cym6tfs+b6v+Eba
mS01ap8Nssbt+NxEXWokDU35JeQNpJK33VQ8NN9MXTCECIT+lrRymoFC7/bHtUbEDngJsBwkKMSQ
7UPo0cngEeu0wAgluEi4uofv7B500QTSL8mF18tYF+fVGIffE2Gu1NbT12UeQHqASiJQfrFf9hgd
/p6ncNqQBZ6Tt+Be3pZUIg/bBItNNqOheuc8H/+EjWSviURx+T6XxvT6yJuJ6WvmjmX5jsOOlVI1
0HeE2l6IZP3+LZLlHRTWDJAWpGUGfb0ipk0JC19o8RRGOTeCE8TQ8W3jN0nwzdDhlPQexATGccZq
CWVWcGxFfmEddcy6NMjhMg9BRQkAmkQxvujhFunVef9TUSBsAv+dEwKbltbC3SiRUNPIfgnoBjdr
ZwXstICKHFqn4sK8dlsrsj6K2lyFxAWz4/hwjhO4fWWjvYaCod1FGx8BO+A8y6cgSxbeUAwOHe3U
hVSUekVi+LEtc5uliyoPDeksDxfIST/3DEv8u1xSN7Stcbaqcw95lcNkyT+tEP0uSpduCT7dLLNM
e9Y4qWKPYfvaeNIEhIembb4MOOuVF0BN5LtWmC4cc2UWbBiOknm4/Iq8nKanVCHNvRRCsx1spHzD
5sdFMZsl1pZU14stqg+hRUaDzUCCjyos4fyUT2abG1QXCQu/USwxpWMVCJNSW2d0A5JrlRc1Ntjy
DonHrCuFdyiFBotxxjKsXlOgB79SLwGLUtYXmvhG8XVw1cw8L+j5XTt6sslMrtMWLkj5jiqwtKDt
oIppyJR0I82LWlIQTR4PO5j+kPaKvxmE3w5hvuMC1AGiLQz2mrZnvpDyy//OehuUGjK1bBvF3h4r
lhO7PrtzCXi+Nq+MXTZePbHlm0vXptiVZ8MZ3xucgdhkwsFx06BY34EjmkMvdid7a8FuBDSdU0jZ
eCuxNFZkG2Mb94D1N1oGiSW8NgleSi/GUZMr5XX2x3B6VMQfKasilwZoiujAJ7xWLaXS1w/dw1mU
HrBTAC7vpN14cnbA3W7ThuCeXPqSVsBPtVgmSFeXzHfa+bQsKBkuN1Y/sRyoQFEq0k776b94/yxI
/44PszP41mjaCs6KB8MV+bi1I0lHgfd5MtXEbAWYjkehHKgbFlHxip2FdRrt+MY74dp/uAlgumwR
EUkRXUw8w4hhrf6hSaxbM4Q324kDXQ08g/enCc36300VCcEUNThJkD41NqnAZAhImUOo9m5Wjfk+
9JaTdyqUSjPI1IGF5mUubcTqTfdwaPGBU98qPGaA1XRgrsUV1m/GAjsrh9ofugN4H6e4qUmDNqFm
YiswfaxP92fbCoTEHAnFQ8PTAw1iC2ZHbaeu3XRR10LrQo8y0nGxPYGdo7abKkPYg16UVxUYFjhL
gHKmaO5CgzFpqr9I40hwDjHztF2GPXgOGpOEWi+gWhkp+CfU+hnnQAwMnQWLuHyjfY3t1ZwzdSLQ
uk3ElDTA63pt5HxiEThOPa1yK9X5xxSEHkrHIAeiQ1wgGrCzmTreimDB6XvDTgBh2sW7dx/7J8g/
u5ed1lb6lq3Bmnock5sy4F3FwVNeJH6rxB8NIaezYqBDOP0BhmF9V2CSEZWVW1aZQwPqvZizcTTy
Bog+iRP1IYF53Y0TxcFwqVO7AKucLcmySAlIcQQ+AXrkVa8Yq3kd4ADHmWkOrqPjvWhQnz3TXzmR
pb5FQTHzwspUxrJJ0TFqw+icDKlyrFaOd7ipQz4OdiTKktTWd9SqFQ8oJEGtcSlFNHCLNpCccZU5
ZYIV9sLVinr6QOjETnJvzPew/+FSfdoA4iJjSrWirDMZxrF7cYMDvK3ctzv78b7b34ilSSUZEa7B
+LryBaJY3BmqVgUEC/UDuWS+uKt4Dup06KxFM5oNAzAfHXxu0SzRNXl6IN6mhUJLz0ncBUuyjWBM
44LOMBFx7pWWmrafiuuUtDGq0lN5seAjwdQFM3jjwXTLqubBhA4cQIF3e9PiN6so9gfFmpcksGYH
1UR1AXO5npddXvDCls505+syUXfJW4htcltAvZ1kVzD1/uPA2Is5Z0M+UPrF3n1vcvJ28b2uO3Ib
eBUHv7xqvebl1H2ekCD3sG7oApHI/heAMISIf899qnjfqgp46+lqsiP5GG+EHAIXpCm4R2FpeYKW
AuwzcauUNOgZFgvuUOHLrJOtbNvNz5ojdb42cf+GWTs8kfcdyoaNrxGwqkIROfJiZzgcrGr71acO
EFKjDMm7lSPHfHk9X61Qiom26Y98nfKyxMPABPOw7edfBUaSo8NdvdoZl4wv0G++iUHjxz+OFr1P
BBqqpZ7UxudflZoeR7c/us25rYrdP5TQyN04D/nGpZzz1GZHPrcpRHWxYS7UxIfpwgmJkfFHyKod
iAtD0R/OCUJfLlqxFeN0XavxWctsTKNxOrxSTxS/KAtwkuruK9ntAc5f5jnjD/JhtRyYlfqmpihB
cqhjdp0zMVy1l4dPzkEjQknLQfvks1b/LrQ0ymKAuAXYyBw1FKnOLqyYNOKRQnnYVtHqpDqOm0Na
RC5iySCjWhiZ+kGMS5RJbu1n/OnLkY7WcNC2JJ45MbUP4G3IRfcLnOaefhsjk5zev0tK9yPsb/H9
sAq5XSluhGz0PxaV5X/m3ux2/2LCOuAeER7BBJ8FLY5n90hB1fKze8w44ub4jahML7s3RffpXQoc
SrU0vnSiRDHeEKUA3G1V9igd0KIEDxdvL4E5VBjnCgscyskd4Rs9Wq26Z1xIBIJ6tDPxjZ6bmC23
mZWD9QrOHrQrFVc0pnLrrzgOv3k3szhajiQqaDq6nhDnvRmfXJODMjFLspyhPTwOv0KhTtFwYsp1
PJ119vJaxq4fXBVdq3oEoIb6ZUcDRJDAOY8JpF9ixq2leT3+rfVz0s3EVe3ZG//WGwHnMDESa+kZ
dQLw5STuHoq+tIQlLnI2yLsKO9ci+6VMxIB6oZTKdtdf6t4d5oiB1kGxQxX425lbJeitxc14wKFE
jmd/p2gz1EdpYt8GwlEU3fiBCUPFAG5fCCOHRALX6TxFC+B+33c5iaqNU8IWF8njMUD2LoWVC++S
ULQWqrl5GqIAgta+kqryjtdL+/WrvifTEe3WjwpFV5VHoI9wbAn1imYn0q+BWawv2rBpkfJ3sH14
vs7WbvPRZYQwx+cQVtcfuRlrigAO932mfJkMhx7rjDINhxKCEHiQ9vm9aZB6etiZAiZyHPMhY8X7
IUc+bO6E0jYMdPvjoAivi9VWxAVQKVJzpYj3LeAQ/jH/guGccJsVaoAf2xLbL+tiV0YL7DXXdm1p
nZcZ463mOu4sLWIkHsZqVzNIUnzHmfoiNTBc2oUJ8tKZeilM3OVEjlK5HxZTfWhkrYfGIKycoBaE
leX0T5eGxtLIkqx47e6CZ/x74OZMQUSSlqqA2leTjc34OEKkl1803ljt5y5vrqqdbm0hiV7dpHXF
5X9zzwNVF/YKZDMP/c/POq2noXsVf8zJKiK8YgRpOFvXOzueU5lGQrFXbXiVanvwPK6Ic/6T3FqF
5XrDXyZXPt+yYwsNToWgVOvZ8qSUQgNl6hnzJvh1h65fopTVp3O680gHl6ilDrrgOGSQ84j/KoIJ
bA/LxULGgoUrwkPPImDiUA58pJQy+90dNvBpAO1NWRkUPqZhYyjGaIneYTqLeZ6VveamNK0wfk9b
Pcg6JzdDSowEWoZ43Rh2jgKcqvUmHVWJ2tfegt4zQFbcA28CWEy//+EPLXDqO0xoPyeeODe7mj8A
TtBLneQcXTyJYdVn8FctsBbKEyen4+M4v0cXYi+5Uf96NfZanVglHlnj1f3W7rsoL6UhkF6mX1qA
RDSTL0Hcj4gKCu+Cm9+jIQB/eGbsdEhAIa1RQHe9iE3+GOl+fr7HvdzIOaqJqCtvJigicpXRiCXX
teDJzgghkphVsP/dHKn9LK38CQGNHIWRSMIw9bGGBzzybtej5xHZO6nmX8ovLYjVNLdJ+mnAZgrp
d8M5OVOsdibarnm/bxlkvss+jc8AgWnPZaTls3Z32fwzrVLTYQu0tT1FfM+iCtNBfDBAAl75d+SG
1hjN+7Uedc7xhLvR9Z1xK+MipEf9hG0yjcP+/jE7BchmqjS01nc/kBDLGN/hTm65Ln5o+krB7rRv
Fl/L94UBISBC5AEWe9lKkrmcwfts6QXF8XcEvTVWsl4MEab5aaFb2dy8l2w9E7mq0O6riIvI37X7
eG7LuwT4t7kNKbCRynoEgXkQrURgtNAksAh9W5iKouAKnoqf4+GBPmKCsRSndUutCEA1W1QowYbI
cTc5CWifRGoq4ITxD1Y7bt1At3crUIqEsZjhkXg3396uOd+c5JHIkx2s9jwNcHotTdy7VRdswGt2
GfvrydXfFpuP+xNyd3AlSjFPNl+/Eu7guz6ndhK4f45P9Qrc9WCwODse0PF78G2P8YglXrv5nU33
8uMNhdOoSd3JVqVgSD4i/5qi1gtZ+2/qYur97WyxpDYW6NzSDuWbtCj94MblRYe8Wfi8w0lPwWv6
44qserOyBeGpR1YXKb65uFV4eDYvMdt1ewjZjWHtBfBHh4/AMHi8wxcMwO5TA5EG1wXIA3MGkYeI
ByzDSvE3xVYoDvMs/koKigpgxobhwyYNsd94go3ThVVDCermMRSppfaU6rZiQsvAGsSCXFiQzHpA
XPsmiopQ/QrEV4AafMqJ9VLdWkidu96yheATC6En+iUg/EeOTYc2SvaU1NV6XkGMmUMFPO58k6Qf
rqA6Z9gWqn//XZ/CEhZg4koTrWpGJIp1qfIjD+WqleQkFnf8MpjYx+jSQmKXy3F2fxJBDDhphKda
3M0DA1BRoX8/uv9c5nSIT2f8yQs0CFhVQFo+Ef5Dy9LZXeHxdzD+JBJ6+PF4mNlmZpUcnPN+Jvz4
aArRSxs4gu/nPSvYzzTepJRhLnQKLT0SH6hl2ekYwiIEM/lLcsg7Okb7FQ4fi/Sg60jJcdnEgIOH
gJ4s4XDPgpdPpzyIzz6Y5FMA7EG3QUi2fE2R5/eKo5kJwxF3QS8Ec3BukaH2X5LJ7pW6m8rtf7Wj
Mls7hSGHecxfuITPufuOetw/sOXkwgosgopQbpE8QjDrO3rMBOoZgFrpvsOaIAoAGW2o8LyPxXGp
/AfjdufSciL/6LBhPoXY8F6GgorahPOfn+tOH9mcQm7WgdHxHiEc7VfU83ZHNCLhSdWMiH+jUiYV
iYTvvQv/FdhJh6WbYqruQ+4F3xlYvXmGcJywA2nRmovGqRS1WLzM2HVYrbrIB8J2fbD1aOjeWCKw
Qz1ki/DRvyDD6hA0FroV9/jHOkutGh/oj6+HggAsvvpgiyOaXvFI7OfkMJRezEAj7rLfOgZy+uvz
mlywvKV+2AnAr9ZqBHsAnhE/EEhqhxzowGkLKryfudwiB9Kp8x0yH6Umg8FLB4Hezh7GLaFNMnH1
Jh7ClUOB/rjHRPEPi1+SAQtCtsrb4mIw5KSqL17d85vboinhZJgRaKTZtyzOIUdX9eZvk/yzt6rc
pNr9/y5ftY+rDoJDVfUn0V29MNouZlcEsVEZrsszfa2/iCJ92rtqZ5ENJK41XaxyqiiXSwUGRE9c
ejTatCSLJOWNPdEzWvvWIlQVtWCxzf5PcaZbToRL+wl2+zjuKxqBAdV0T7RYPJuP/L9bAknPQyDc
JlQo0itTR6QvVA5P8Awh845gdE6CxABlq+Ccg+B1/jYxnCNQffVrnKkD21BISAqKrFLTmF2duVjv
aL2tPs9Jv/ZiqeoCQn+wIjdnwiiAcVeNmXB2ytETeeywZv9vUaNHH0x+kpaDR7MW3TkQx41jbu3u
kG9Jt+oWCPUr+3KPOobwDTBUgYQcK/GkzSuhLNjiwAGQE4BWZ2gUve/YbdQEakQrHtRRhHdOkiKf
+BYzeouXBOD3I/GtsiS2FSXHN0tMdW92iQn+s5ThO/Pw95IO3MOXm6D5J0VeXtlw49QW3sPJSbCL
UYnacgaVIaUIGHikXynccslEJrru6Sk40GmQ4GdkVKS7GYBQ8c5/Dh/heE4Xa75YQ1qxggCACp+P
Z2Zez7cYlEz/7SLYjVo5eU5/ci5lvL+mVovtPG2MJJf5odKNNJzVTjHOhX8jDcOcHcmdy3+4INP4
2O+7/xJZRVH82xy+D9KCgzKKFB2hJhQkjz0FKUxwaA7qvjXMGtjcSZ13T2xr7hLzwqc6Ss4Ovd+/
vQt7n7oZLpV66HZJAc0zzOAzvb3gyFHzIvztT7zC+rePlmNwyh5Tnk1cPDdrAhLVIyW4JdztiKj5
Rqguv859jnGcNkblf9RX/OZ+Pr3WPWpLjh0fnNrkeXeIjK+ZGPuaMmMrHPvhKfHhWmDVjGEeQOxa
tyAqOwdNr7O6xGzUUX5B2BOP6i80eh7E9Hgqp5I/6XiJBDA0VOK+AzPdrU0dRHcizeaFovdVQMgw
lIGP2Mu+eYbv5zkLkkaGN5osuiSlxLICWzR1dnrrGHgIpCTp1fXx0mgXTQV18s9cRLAAPofgjHDM
nZW5MENUt9FnjnuxRXvA5xB+VhTYeF/AXqzkCuJOYPpyDi0Hbv0TOBCH2sNSorbgaacuMijkr57t
v5aEU3QSOSbFb752mKCEx3MeLxxmf0/kQ4zNSbO0Dcz1vojKMNs1k7ZvW+cK0ksj2DTIX9duyvnR
9KjLBWMsgMrkBKVJDZKyygJzETRpjxO80Y5tpsUScwp9aAGB8hy8yxrsB5J4R47TrGMhXIxCQWGx
s9qp4fTm0zjb/uFRKLS/uIEU67Vh+T/LBsKAzqcLZVHOnbhNmjYowMzpAjTxpXcWWP2AvomLIclL
PP4aLL3bgv32cL2CBSmiEVYj+yYFgx/6Lqg0d5TwAddIvsu2tGUv5heWsot40jVmg92AkoljmNuX
I8cO0p6idQ5xQ9tfBrQLx/BYbGFPLHSXnnvOxdQoY7BX+OYg2YHE2RlaGZHWqIBPOg1qMmywKloG
TeTJhCNUhm5y/HFa81bi5JRh6qshx9BScXXha+OeRR+20buu5Jy2FVhRIVBnA95GrnT2gG3Psp7z
4gjiCkJ9m0ZlOTDYf5neV6vAUR5K8rCl6GSjJV15THEiS7CIAYABzJ7IBudJjPEPRcPUjdCu4BYp
RP/W1cfDU5McmP2wL6zpI9ZAt9F9/O35JjTiNb74FyA26Bm6CUPIBVfCmOpYs5oHi83Z0NVb1s2A
vW1rajLvVSP+/YkoVnOfufgTEqlw63TwMcHdM49SrQdbLUbp98h6kZLM8UZbZmUjfc/z5TJFepVb
k979CPwoskNqs6F60bE2tPKyDyyPAe2J3Wvlq3UfwalMq4i9ZP2AbGSbUPcXFiOs2y4kEwSTt0uP
e3E3V06syKS4X/VFSb2m0BtfdQrvyhP7cfIP7CJAdkM/vhmal6UBFyulBq3n1UD7YKPD1pfAR8V2
NhJRIa9JB3RAiJ4fxt6VwvttMFrNYoUIQrY7ziCoyJSWYrMkYtbsUd+i+ByXyTIPp4k6IWmg6BUv
EsQQhQzwvo+gJ7vKwlOLfUj5spldP2TH49Ba6ktVVYx+7ogZgkYtU1f9ex0G2uvpD06MPChMbsG2
cJmcbQQbiWUC8BLqT80iYlQebvNClQ3j+d79ZhGY04dUp5ZWcNTB2UKgZ7dJnx4EtEe6EzqxCjtQ
dpqQdcmUDER5fMLuY7Lkgh4sH708vQFT2U3ZtFiXTfnUKBHkOUNjSozU8MXXctjeQlAbOd6gOy1M
oF2M0mSwyrgQr56x9aM974yC2py/ZhbOK6qwcCVaMlN1XxFJTy/yomZMeJsxRA71mcoTYSjO3K2V
OpkctJjdLDC0gYK5SwZKDkhfIX2pyYl/oG2ajU92O/+Y6oatndS7jhZhPWki+ezk0J3asvo5PVDe
EhUGteACXmIJ9cgBjoJiaLmsJdEYWdLQKCC8zctx83XCC/x2Xdm7rcji2m8jQFkvS4GOW5ddc+nM
IGfnb/Jww9YHgghDiTlmpw17HBlsulp8U3fkHTCHibN7lqzxxaOPX+QiA7WWni4iKHt8Pz6/rrcl
X78I5eVZV+bvMRHTeHUBTzbTAe1Q6s6pZxb5ColT9SuPTmivLN3EpIk9FDY93WikW0USqu9U4FbT
kIduQIrF4Fk54cQEu/3yJUUe6e5Ji087lzLHTisHGoy7Neg2DYl1AQl/5oclbfsqvrTfKyi6RQT4
dqepk+avU5Bw1/oESZWFtm6pTRLY3+UjKkyxsuSd8RPb9t7Pzngkt8V7O5gASuQ7tiD/MFrWVyTn
nQpUrnxXg9x6j5iCudf9HcPDwAoYT+3Zp4Yv3+t36Hnr76eWAFObq2aG7HnNQXWuTSv/nz+4zbmn
Ol2agdcfyghfkTM05xTd8SQ3ia5kJY7T1TEr9IcXQC4o5v1uWPVQLkkxiSgmj7euHGMEYNJNsLZn
2JX6qd3PamIZnHFL3Gs2GOmYeBh2NV+ViGqRvnp0YrwvlOzNTHnOxccoYzfFT5Frx8JuXr5RZ+Fc
I8g205evBAMkqWAJbRnrqupN0PByNjqkhE6O93RUJXA4HHrNiy1gdaCl+3nIV510Ci0N0l1jrOwW
6Rc3IRcveS9fcrcYr4Tb1EOw4ctC0h01ROitrLU2ThacJ48xuYdEaJ69azjvpYidXRf+iXPG/X7p
D5ORu8TJQYSEN38peUKZQrr28vGPWCIlS3/yvjKGBmJsCdzkSooM+t41mY4M5YHDAVwiebgbYaEk
tjZlOuMEzbzBD8bPI1u++H8R/ArX4Qrj2BuVtAcnvBEWdKfEV4vZDK80t8A8NaexJGs6QvrxThWi
dFCIm0h5wpo1A14NlrI9kwXhyUIIybVCrcuTYfhKbwJxI7RBCtsu1yq1u3tlDi385BRIEfa5Fy7W
8+viT6IN/Fd3He7Y8J/8Odg9ILHdeUMGsmhT3TCpoaXIx+Odcgvm4d5rzPlAdEvT7cPyIa/DVe6e
9xSHCRMO/5we/rRhVvW4GY1z2HpcQrF8gJWziNDRgrR+tweu+oZhyiwfyHT5/1qIeYBVhtE4mICU
ZRWrsCMOLB2w+fdq9AJi4tx95NsRSCnKlGEyQBXaIN7DJU3r4QL1onUeNFz+aXGV2KIqo+/EBwB0
kyuGzW+uX/BJ6UC7uButw22gzFKX8PVZHZYUiqbjdKCPoEHwQtBgks+iXS6FW8UIcKYlhsitk9Sp
Q2u3f/Zwe1UYOli8qFV1vhxw/2dKvMwbNY+8LPx3eyEfiQO1cqwowHFJgiBEd0DBV0zZJkYCWs0r
E8U5LYR+OclvNH/mgpafT8FGGhrUAPOvpFsPY8KLZ/J2wL1477yjY7ud4Zgv6pI5MgQfFn05YbpG
qnv0CqX9gccV5CJ/rE3lT5I7BJ0RB8dcpHAv2futW1fdNmE+RFuH68yljX3jNkvO06EUXXiwEm7m
Aq6FpJVKcCdHipxNSuQPDLfxouuhZgQM/3JbtLRH2YHU16iRgA8+9Kgron0+EyYmXT0jn4r6j7kQ
XtFBh9TU3Pzs4glJtrp93CeQoAkj4iKJanTCwWv6SiasTU6tTW+t1tqdJvgtsfi+sVmYn3L8MOGq
5D9I4YAKJS3G8Ymkn03LhIZ/MTYeI9QNrVgqGR1S9AXS8li2TqtxsW1ZcBbYhiCCTwngdxjUYMrF
aeGfcM0icEcNoZJaMuEzdH9c2nkdlTdm0bgkrRlffdCwdnHHdjaPccRaETbYAbeecVGnFCEsxHBj
kKLFpdgYq7f07qFKiX9kL+Vwffkiuma4YE0Ll26i7oesaHUAWJpW7NS97SHBpqRpWpT/6gbR09lh
Ra1nClBe+eD0go4TckJI3j4zXxClC3Ie8a5WtBSDurvoPiixP/8xHsV4eTUguv/zl5MeMtOFj7Nb
3JhidCbxdryKNHuSRBZ1eKEpgmXOe52tYlanPtdiySfgVwWkUovIr80Kki5mKrOBV5Yo+QgFLikm
+wqFdorf/TyYEwR+QwFmdVFDP6AJDA/YxkqJ59He7gvetMvgnNHEmwGID/nLUa2w3G6jUeAuKOZC
FGvXNK/W5h+N3tG/ysFOJ28GQzjmX/8tBBj2DWEfHLz5A9alP/lgnRwVm1HKOlzz6tt4EE7Vo/M4
CyCCUhIEWf8Tqfn/Cl41fL00gWcJCTjLkWb7pqHzNduw5sw+4dqBc11W9Lmz341L69bEdR4o977Z
GO921fPDaePyv5oaUaPd0LaR/Fzkb+NyI5Dj215/9i08I38QXVTgmc+mjmLbwq9zHHEj61G/1E+Q
xWZTho34T76OZadvYrKRX2ZQhOUpLb8Lcveey+F2CEFq3E37PCkmGPbCpGj4fmsUlS73yxwfxgRl
e27ta7FYeII+j4/wVCiNgfmoa9ArIeefp/bQtSZuT4LeNpXjTdYb+CmBnoqYBdWtmQnpZTXvLoc6
WT/MwBW3KKLHInHmF2S4qdY/bo1LF/RNIY89t73f+Qfs6fHL3nLIuddFzb1e7RHwXC+X5RYa5oZ+
rPrxJ85Z4z7DPwf/xoPeadIh8WGXCWGgiWP3PCel76EZ2NAo+cXC1lnLQuEvoWgsF6gpkQH3R9w5
yQfWotOnYjUo68yil1IPbvmqfOnUd/gp7BYW6nExdCuya5QFGRcZU1nypyHEaA5K6qERiKinQmCO
jCXeW0nyhseRt+IkTdamZjIJl/La6uw94yGXdoqecjjGCArEA3BeOj0VfDqRGfbDFpcv/Gkjlc/P
RFGI50xQ1nB4T1m8fdUlwynAe9K6l66En+/8YGY1djMsMsU2ApLdJyj3qv/66qqPn937SFcEzHdy
zN6v3c0yFBeAKsQy+RoJHm9Tod8hK5rQ6rgdy2wj2Q5R3WkfRpTjFOKYnDRQeDt+QQXIkSkOslOh
7wU0OupemCvR7o5NfVic83IK5CEDD2WFXO2PF1XryD/lSqqNoHqhnEq4l3CRZEDi6gi2vKeUJVKv
Iym6eQGZO4hUtiES5ka5a42Or9Xv+l7mjyJ467lXNJiWUjOu5uYT1Dz8K0E2b4DJNsTo8ac0PZ0m
VSaWTaY2MJj+pntZUyIoeg4e6exIKvIIVv4BIHSN56AAFWlnuhTN35iuY0Bt6FLnZ9FlqCXcqnzc
JjU/L6/o6NKCcYq5V6wZuc7fHJVubAHZ7O9JmLliaYT1WVgBzLPg4USJz5qi/uu65E6G/S/CR6ec
eg7tFsaP8HLU3/r7Kg4cglfozIUW5ouLUEL+bNhLv2CMCgJThbgFsW8w8XPqiWinRkCoKmsc6hgT
0q72chzXx21BwWHPfKBcyWas9yoWIpdJqxvjaio1BO2v0hfD9FRSS8N7c8dak4jyjFJEC1DVtoX3
6suP4BIbint+a/cY6vFUpxw0gd/ay6SZK39GNvnhoTB/JE9oDFLdj1TYZ+sM1UuGNEfOU33yRfL6
sJ1xzZBwOMRCJIAUOYV9y2Mp1qaST9xJtXkJZ7qAdUN8dsVOuG/G1xBfY9pxjtlnFTEn0dc+salv
USdKDnOrXDwea6NDo2Zq9yvP5eeAv2hL2SQrdoMudzcR0i3Ukt9aoUvZzysa3Ucw17+2PvFPGXk+
9FSgD9bLJnmPbxCvi3727j97a7b4cNYBsNXyBivm3eo9x+9uhh+hljyhKcwIX+ZOiIuaZvnisRKL
a8V5ZIR3vy/LDE+CVgNzOuztYF51N2/+eeKtM5ryljSebVCAxkF6kMuibH1g0EbItKEpOGIKACmd
5bfBYg3HzVPmiTEfprctgCGOCISOEERDK6mxm1jMkMNrqJ5YU+sLl4JTxR02zUipfm6Sp/GTv8/9
gQzujg8ymkwprd+x8hotj3CSK+SmGJ6pGlLNh628tYFDIufyLsYne6XEg9q6TiBH+CBpHQM96wiu
2/QZIheMRQKmZh0dXEhg80XvDDWE42lQ1BpvkgsFVvFcBPVtMAZg/bI2C5d/4Dwz+DTgo0qB57wV
/FC4Wg1HcAXWAa9ywEb/kSKoSGuny0xH/APcjSg7IrtArNZpKJFoPPpDyH7bJjJBjKgbw0Bgug+z
jzZolSjuGpxqpZZ3ko/YAfHVH0jIaf0l0CYd1LJn+COQl6bAp4hEJoJszWvwPKtl5wTzFvU3+m+e
pi1w1iMCAvXYpnhGtXSZtUSEdEtmCbuoWpoWFVFvp1paoO+D5+mLz6+KcUjO2M1zL833pFy8WYQ0
eYE1EI8G3D+2VlKkNNxH3NI/qm3UHknUxvWbVqMUDvcTdF7q1q1e74uYkeXJggMmKaV2GiYCD4sm
9gE1tMbWs9prqnfPnc5izsPETW/4h4PqV86ZcrlKEDB2Sq/aRf4uUPnWn2EYDjZjvZfQssLGdt+q
+27d/qQcux6BUR9E5Bl+LV+syhC0lj9NPNsUw891vRLoMvJBSv0jZjyNK4TFMEDToKPGrBxka4Fu
HUGAR5EP/231qCB/FS1M0aKwEl1XXn8VMlf214pQIaaQq23wNdFTClrOyq4KmMTCsnQG+G4NHKYx
BEK2Eai3M23EPLEl9cbxdQm6nHbTj9p/zuuW3LhzG+I9BExzqkmfTTeOjBSvfJv/KlBhMYbXNcqC
OtWzw/kivqdDvQIsONnFoNA4RGeXNXMIlNktH8yI5BW6zcM9Z06pdMC9W4XOzguKCmgsw2XOyAms
FKdISIhkGnh/oKnVWyzt7ar+bBTIIGRVozX63YzMuGvCg60E2RNIW5numfQaAQj73mFo3+Gxi5bR
o2mOXqWyP/nmWslf/GmV7Fltq0bmlG+zhsq52qx+xOhmvg22TT6lHecq/yZSSBh7qmKxaDuY9u0l
PgW0XVJVPkcKJmZKt57EzDTYd7srt+vgHpQxkcJcYothtwB+/XNRRryfqwOsHd8dxI9mt8S6tVng
DK2BCsIZUPSpjvicIYrtcze798sJJUsKk0Pad2WEB07xM+PclCUxsRwA4Zx1ugOF6RbF2BV7mDpX
8dBRxG91igGw5rcyDP+aJyurHqgNeiiK8R+VPTyW3dVVHwTMNlM5qagtqHjpnhapFfzvFSR1Pc91
Nw3HJYIIneE4miG1xl288RFJ1G2mR36lM2wMGx2vdDVULIEbieiRc76Pw+ptH5B+5ZPlwddBXpMV
xo9Bu3+mSD/OCOD+AZmDRgAdhF7MfpLID2EU2aLK++leUBllkYh1vy6y0niMpKI4v3w2P3CN5UQp
BbRvjWhJt+PLsZEX3F5Lb9mqFWyeSgHt3tKT6J/FpE/Y3bvjpCkcDQRl7USLgT1hNGdPGBDqogbL
UuGJ0QCyyvIMdID/Tonn84t7Ty3sqtvCm9Gb01EAQhKYoln4XcytleE6cpelB6FnNTkyCjy8H4c3
AmQGptxAg0X2DxGXDf0HNbGhtuLSU7R+0ZO4a5YoOYggweA58z5UhdOYwsCf4yGARFsVg4KyxtAS
TgO4XV9aYaHDssKDoe6eSbleVCvbYIhrVInMwyJbRztdgXTmWvWQCaYREqG4s7uAD5ZZIJnm2qgq
CBUuQkpX//4VjGqkTmieJiX7OYz6b5oHWzSRScKAgGCSfRRVV2T/+NfQ08AXDpU9uCHqLbP1Xz2h
x9SFRnmdXDs316MJI++JgOxnrAUiRyIKhH3oeYdgNZ7PdQ5dX5fpa2LKLgVQJedNSKbO+2JZOmg5
kkSpUBgD36LF7YzRA5j6rjfgRBOTiIXlLQMc6kxZH30R96CUUoCTZg6s7BrXKup3GGSNXxxcH07o
DXtolR4MluAwKxXqKBcq0ZNpln9UEEz59HREo+KS72QjU0Xdtq8K53DOwOrKPClw4zml5mC916DF
yLNSv8UBylAczXgiPOjWNpLoBuJ7rp3njnQrvC5FNP5paHOwL+HxZ/G0UAVhvScc3kArGz3sLNlA
dt24DHSXt/3v/4h9XBSKPfube1s+rtzufr0to/XXWcXrzAZmO4iPbk1cHdsrMcGEg39liWy8PAy1
/sxn1dWwm1iQignLxeBtmzK/rte/mZByPqJVNQ8cNFvY8JfCGmdVAsUpbVmO2NROPlP5nyaOtgJM
1ccrAffnXRVpwRsCU8bPV07eR534mZQazrrsyn2vKED4MApdxZ1gpYvV4zgOQTtQRW/lpByN1pYV
QBOMOduNABI9qH+r4Rc6W73kheh8+p8O/RIqljiqlzPoDFW+l1cAbXVnQg6NZBsX0vLZ3w79bMOL
1jQyJi9TPzpDrMSVqUZgbs3NtvKXSDZWvOm2Tx0Ga0i7UR0EEjaI5HjSTWhavyy/82T0qRYUhy6Y
WY0TJNXppio6DkTXeyCagG0pQi97HX5bJZqH07KziGfCyX8cGAq/uHHJfQOYYCSzmQUX0L2XxWZo
bXVdmJnX7JR3ms2UYMoeiXUgGjvsoH79fhzZ4Q9IxwemAJ8al7cYvPBs+Xyh8+efl8sDSBhHWyHQ
gsqFgaFvQF1Yfl11vSh1QumuyugS6eT+/k3ieDznrD90bPJZARyGJ6zGeWjHVQxOpHnexkicUCUz
zoyM8e3wP3mpYvXK9ECAGTGHFxod1w0atvRClx8Wd1thnbPW8stQinI5OptKpHPK8XgFTuiNNMMf
jhh6VMhab01ZaigpFa6/L3m4gnfVw87eEOju9KXc/M33SvghX008nOmFBdl+Ts/boHistJwh0ZUD
TFLworb5jV7FeBe6MNGYGNOA+Hp83IF7yjzVlgBewZBA/1OA3FeXto5REhRlDLQqElRG4E7NE1CB
w1LY3wLdAL3q8V7ov4qRbxTA3Z7z+7V00F67r+BynCrUh/jIsryMLLXy7MKa/YCb+e/ek+UgAuZJ
jsQaBysQCQQMkWysoKvmN36KH+NcoOCwIKakWiyG8rgn6msyZ3rnm+vTejrgyuStoKSxRHaWUqrv
ZWNXz2KDhZVTvBPvhOxmJc/chcvYzcBHEukdrvfAjTsJMM2/xGhdKxhMkL/CYHPS5uspLvgwAwzL
aiW3avrXBSPDfHI98FSf3rkkq9NzXF09YNJn0C9rJra5u0tEmvDOmTlG9QioQMTXD4Lpwmfa2dgP
Rumsa6fcUO9X/yeWgacx1KKerRLdi3GvtujizLITHbMtUaVMgWP1sI74S2Y8hoM/oMa+/eO404eV
n3/Jv8iFKU4zqaf3PuypKNq6Y4XEFYdA93ZxbmkKJGdhT3SlhxHfnFgkx5t3+lJAuD87kL8qbTlV
A51FAcQZ1jjolpWpXIV0JVUvx9b+5WtmqGyFuVF/O7vaBH33xZknXzzUPSCIqYNwsxPPJfovqyv9
sF/0a7sbh6tqP34beIgUlK1elg4k38yjhmatP9lsafXI0mNMjzgk2RjJkXlxeS3cSj3mY5c1VYQq
68aSKbQnp1paOD4nw8ghiJ+nvx9xcfA4fri732fAXYuCL1QvsPudMRhtzIqtXDtY3Tng5JTd8NVv
HPRy78gyKgvRiB6D5ANrX/Sr14CJUDTIIzhJuyBdNTpdOa2cy78UJGL54DkotPum6xaxKwe0BZ6B
SRcWjOldK2A/ULHg0WBx083R3UQ4llI8JvKG3yetUol50SsN2xBWJTNaFWCNFa4x6DS3OU6ssBCE
t9w42ud36uXiworx7jlKXkXKGaVi8kKaTim0K48++OXTvSSTJFXGbAak/1/mfUNmlZlSFi9v0IQm
/Iars9D9Je32G/Z/6XtOwS/wl3G8r/LbkwswNSbJ+FXwHOcwjgSqadgzuxmlFI+RsZhXMWyYgMKy
7sXcmAHig3jMJmvv5jD8G0gmRS+R6q0TuReAoKNA91xvr0Pi/BTY1GynONbnIZho786dcr2bW+ud
F9H+/xag42NRIAP39hZvnA+sTvnhoWiFyPTe2V2APvoMeKzkkMMSDYj7JRfZq5mnGgmxuRqKKMgf
z0c9uqxMwq9rK2LuBeouuqyPaSRN+rkjnYWIc73K/zSGxLYeGtMjBXHjl6n5riiEGO5PW66VMK1L
4CGiyYbOpkqFC/vdh+k5+Qi91Fwg7txo2HriFbxbMKSg59a3HozUKrI4LZB2eaA+t8sWid2z21n+
HPBOoCiI+KUt/sANMpPA49LXMmg3uGp20wlVgpScG1Rh/JImpzpK3KSlN59V19DeaLzMVbkNuDRU
vyADV75mqr7pO34G6yF0PyOeKXdngMrE0KNvFmnbdMstcgnXhtx7U+6UMFtYP1Ay3Ge3qICSFuZe
oAoKwgtriDItTYiOcBQTcrY82MoTeXKLOYRK7+HGriQL4xwk0b0PivLjqX0PWEFUvMx5XmRd/8Ea
l7Qhu+kvqbBW1cyOB4ltJ1mv2v88L2LeKpvV/6WrgYD+wFD923GYf/0G5q3yHPwT1v2SnA8HOj0t
7f93yM3wtgFKEHD3ENbeByWiSmgO/iW+09DV0ZNXbcL1KOQg/wQwHdEMZfs87ArSaRqMpjMbiWSa
2m2eyIdXYBYIf3ZkgD9dffZ4ZJvYQ4yIHuzV0yDShLVgQF8Jvhwu6bzhigEoa+UTXEJJpImsZIRp
27FNlY5yyBOGkTK4J7IzZ7+/tjVi/wbbek1FFpkwowUw+P29AON7P05WTHvoAK3YL/zzdtv0D2Pe
XyxrnpGtKcsDZqvIuiG+7nFEdlv/6WCl/P+6e22WUhm+jwRtXJIxG8XLA5SpBymifF9vOmg/VtUf
g/p0XLz4kfXYZfntaE7mxwPmy+f9AIMN81y87bPw7B2x5UCZLnS2mMRFrysLk10Zmb+0KS9nj0GE
riqZDB1K+5W2Cd1qtGYXZvCWoEt4j3+mUh03xcA0r2zdyZ2FZKYYYI6C1w+443nW/Ib+tQetm3pH
2rzQukpcRnoypwjSiu0W0ZPsp1REdVkUQYvul9Ty/mAbeQ/w96xHr8gPKridSLcRFu+HDhlCYjAO
eX241Zgrd85+jWc5iTfdmyezYN+m7rfXQgjcjNCR/3zRtIwtjoOP9z3VZVvuTuiE5g4Nc/I6LmHY
KI/B03BcZDc7zPCxoi86Lzs0PEYtw36Ev+3bY/68lWl3F3TDApEKGiUTNaQblVoWRnakoYm/W7lP
OEYwjM6DCBuaU+XXGR5LvVX5coxHswHFmML8BE7wZ7dOrQ66KHgwa8MxMcqFUuleoKpZNrqhFUq2
diGvi6ckrdjQirlN0qo3LWwto9DbuZZYstyRsJt9geA44XU3XuDC6TJPBMjQ5ZjJvEEcFR2Kda3R
FCr3d50aRL2C4nutdO0v0V27ER0hbzh8RSw1JOuofXdswftmxFa4bVaXxtpwgl/SctcGriIlKmNQ
srm0a7OFk2W2gyamo1HFJVrphW2CuAhjvftKLT6N3ChX303kPmqCizgriJaCIW5eryMKqKzdZwRO
h9P3RZ+D13fwwhzDQo1kAYYx0Od9xI45JzuDj0rBbvmPPpTiUuH02RqZWrD3XOEGvbaHNa7tvGoN
Y8JLYEieMiplAHw+7PvU3N0S3qP3L3GyIdnwlDpXRsIfgIIvyUuJcKiY7RJBmOKwXG0mOPvGxYeL
WnOcpM3xyhkRrQm7A+YRDXMUcL08aK7m9a3zNx2fQN2oEiJX159PYhO/J1K6/htokRMlOq13ElkM
kdBle3Jzt1YVgu+7Xdtgu3A0h1AZUoTCnLrZE4b3/peaE0/QjvhXOeuMyPnbS9JIWFU+ngFLomKB
Wxr3paPz/1VREFE6Z5jUj+wtq2t1DAOjqga7E7goNsrDPQzYDaG2oA8ktgfCTKjgE9mFTsWNnsIm
dYd4eyLkjyHy1hG5wvIXJq9GMifwwFKALnD9IcBieYuAeYdamYeq69V+8sVc1uXznjkh3SRONe4Z
ZSVDI9jIhMg0zGU6LwoqYlu30inIWAK/PwJa6aQmfLee8qR8V2EdtgusFo6Norucg1QC1rFzgwr7
QSPZXlbS9Ni9WmJW7KDAB9id36fpe4Hvas5veFdbAe8ME852ywdPFCIVQS7HeZPrnFMrLioXC8xV
p+FCBCHj6cQ4Et0q69U+ygEfzVvj5QDIhL8TV2cqc3PGcyocvk25I1SAGGPtFFFn5Bc2+wgXqr+f
zVqNBMf0V1QR4Kp5nOM7Mr9vffGkhaNU/5/w14vsS+LJw5ANes/UOl1o9Lz5cgFs8mMl0UY/B9Rv
jSXm1uXVsCp4XDSnSpyuw/SxRgcWPZQgEoV0j0IMystqQrNL29TuqnHtvxU803Mo4hIBMz5ywlFW
NGW1t9iH4TJcuYRpSLDsBc6gXytEOXFE/M3/gsqsS1D6bAPTMUKEoPPd1OJu1bkbUjkXxIu2lJ9r
UIiw4YfhIDnSbYnkLiA3Q/e72PzQVAwCu2OFH/K94dsGV7g+GDp2/Tdgj//TjIIr2EEtbmGuBTdK
mMQ7gW0CCeTJLTgjIuK7a30HxrYSxE5ZYs0O4sgm6d5orGDIzweXXbswP+bu5LGZrgChNrZ4k3dU
TTDj0T2dOFAFfNJ4dBnd8Ww30wcniNUBS+XYEzw/VKM1QNszPCEQQrxusLdj8ewTe8QG4hjKjWOD
9rqISr3HZAfM8RMWxuwqn4XXtwmE6wZ64RiU98Z1SWj7AOoXiQ+DHqmWF/N0QjTD9o3MXXaMgDyT
2YNNL/M1lv7BJflUZBZfCV5uSCyaWsV9NomiyfeFkkfL0EBWG20KDkUR34bg2fdKYmk+Nri6WQeU
gobmN5FLf5CKcVYVMmGPnFFdh5hgmVXX2KnQhhvqixP7/fG5VRnXRSyLttVkAlTCDQtsSs3QpAZO
duJMkat73bWHc06Pslk97sxtKvaMjCGmiF9AGZsReijUuj1IZ0xruinzzP+RxPW+jgnkvb3eav05
3R/KplZkln11kpjRfIvDstqeHtRjRcs+nt3XhpBMsO8c50dXhi58oHSB83PPsBO/tI8FL5Rm6NGB
11OKvSyWkt1fFBp9vdG9FGSjHRBcJme6KFfqTB1ApTn/fEUojby2Xu0q0RCX3qeYQ4I5pyjrBO51
wpAkeCuDCynw97G4kZBt23YOgecRtgQRZh4VB2mAEY4GB9nynAQAuNT6zlesuWvAvRIbC4lNAQkI
JSdEUDYm5lqHH9/i/SPqnZ1YKnmXduhNblgUbf8rMmBOMHLvK/0xscZbXKJS5ZbboM5hm/WbgmyW
1Yuor32fUKCh5gOsxC8JPuwAk5G2e/gREM6FiRE37BUCRySzKZW21S1xyXybApmnVR5vsHThR0A9
nzjGJzvUbtx0PPnprpLKlNrICClHRk2gaOxAkHsU2yliQSjdGApJiAKBYV5UlZEnVND5KUOx16O+
EeGwqg6KdIaq0iSCq7F5A2lQbBddOao5kBJJC1suXQGuofICoRWLoHOuxk6xP4/DRdbXDharpuJj
klON8HYgbTZB4w64kn9QMLnvq3QTI8jBT1mgO/P2m5vfAg7WPi2cS/NRfBnPiRXCNVK2yRnEW19F
CtPrEWxWJVsl7TFv+0A4bVj97ssbqB0RZqb5mbrb/DpeS6BCWRs5lkKBGDUnQ70foJtKQcXYcsmo
pEl5qtgCx9ZnKjj6Gnf9LK0iG+LYunU0Q7hOoEs3FQNkIPZceSOAgiEHaiAfYgZeSu7TQ4yumBXC
ymcKVIWymFZHgSAxGkDMBTOho15Jbq7YwM9V50pKkJMU+5njlgV8zHbxWHi7Fo2/iKNkA/zsHfu7
c7GZV/PgmqW19X4KlqyBqWKfDU6GeJdePEeDbPPPecbuau5LXL5uQ8Fv2XRqo0LEmByuNWpfRLub
JLdchNnJW6FEywF96+U6WHW7ZfkIK1J2aCcDxstbs73NUr61PFp0kGAuwesv1zwm0D6k5YPaNXQT
yQeC5GNgwRQEfxMh3UVrRXF6LSDNWlmWrUGzsrr5Qr7c9eM5xv3DAuwsioAQ0W2qH3WwsD9bccbE
XgXNGdqat/J91H+D/+AUc+8ahIl7TL4Ec5uevMGHcY8eUyOxsHVq87uPzLNWE3VHZKYJ+7wXM/eQ
kOAhWX4iqg3R/ujyPXFik2sDsKMv8DeVWzmtM/XBUJpKVMxRRocIrqH/1Mo0gnQadtMOuJte6gbs
4B+9aCoWQNN3sONQztNWjxpT615LhOCiLhFjye/Uze/NkulUqtgxwb7f3aLG0m8NG4PRXWIgksax
IMBazwFxSlhGhIk+d2uNQmj18+fAHRPfuit8Sr174hZuB504rVTsxAt3fAov7oUP9jNCdh2N6nxU
b8LHssy5M0ei/+YU81YQPSgw3kT1c3iblR8cfMaWsbXeIlOG8JOe/xExolMVmpYryijkcTlmR7vd
IyBYKNBr5g30Tg2wgC3ZnIPS82JmQBSjogd68PLatQ1Ts/arM8mjv4GNciQIV4zNWo/ZtgwVNV8d
2652ovrbNgpjllolfjCglS3Tqts02UzfIZBvYGh4Na+VaAUSsJhaxtS1y8vZ4TkKTHr9og0rXUay
0xriOfZD0Id6bId+umUaQt3ouqa+TuJkaHFCfIdhyIn1I6qBzGuR57TC/1Syvtn2We2FiCOdmoiH
vNj+UaYtUe2cHpTbHR+XhWd+1zNrRoaG3+8oWVTqHD7Ksh2mCE7n4XTieTKsmpZcu7mzJFk9rhRH
aAWm0kG4Ksabs/AslHKANRspcSQjzSzXHJd7wXQxsNnPdJnbcgUEekMHkRdOH2oWZ+GnPcBMBbG9
WgdNsLsXoWY0sSUpQv2Uqp0cPXUuHPvOTIdHPB1kgaiG8Wf7Q1E3OBMuulQb+/RPhpwu84zW9G3g
Cy9TdgL898gKmr3FRmcXgZW3vwALJf9gN6mkYS+xIQ0vlW5dJqeDlyX211Qz+GCkBrMNpGkyzDdQ
eUo+PGtzrOxepwir22/RxEOJm69XChDmggO6mDGQZc1BoscgkK0qlbh6eRq7AxfGSzA1Y+mQ4c5F
5dsOO94ggt5JMdTClTfRIiwm5iLbxc4U33m6/E0gGPgPYW6LZJhMbtNwWcJlD49vjfCmqiwhq1jY
xtHpbl6jZClqkB0pqO7Y8PR3t+68fbpbVvAY0ODMiVKNKQPgZ7vjXLSokqZeNG9bN7MqSOnqgqwz
ej0xG4nyLOQanBgEtrVHb2aAmcDtVgkDdBQeuVP+/hWGzUI5AjDqAoQbMcV4g6OAjh8ibqON99L4
S+Cmge8Lehoj4x1aQjgm/PAvVVovh6h97YwdnTz9/kqdsQzemqR3DpOirkxQJRC+3lfP1BdK6XcO
dblT+etslFztrBuHxCLG0YM7FALF3QQHObleMSolQODLqyJ7rw7eQrzHxtosZ/6p7Uz1Oav79nWa
LLdQIuxfUz8ufe2nJHQ0Q/ek/XyWl71G0po1QNYPj6LFOCSKQ0WFCxU1usGToAnxkReDAbCC5mbv
nvcFzdz40fBhoHkpHJYf+KTf9zT1zRFQtSPnuaw6IEVeD/5+pK57pguNZcJmREUNe1T2N+DZpaJC
iK0665WjXwsvNqd43xDV1oeMdkOyc9qA6gTFZUBS71kBD/VWO5aBqWUkhyL51xabhvrD40jDswYn
BXCSQl5xWUwmzpx65DjrrZmiFIkkBtpr9TMPMm8GkMy8332ycX8SrwwNE9dD/nU/9iwXc/4rahvj
mrodHLeuzCncfp0xobYjmZeXD1z90lcJhBcpUERskyDMfKFiFBzPQ8ydPPJKvR+F92ZLqH0e+E0e
3vHvIKLkTlbnaWW8C16NjpRdY+fM14yHrT11aBnNQlbOODlMAFqDms2Mql54C3yIEcGSgcxXpDGT
6c+5T/N0AkoqweJA13hNwaYAANfWXSy4xx737LFNCaowvpfwjaDZmIJ1HDtkYzn9stCGxG5CPjZ0
ocYWEGkVlpqBFHYJg+tD+Rv9ItsNY2rC8q7efTvmuPsuoA37r21lp8etSjfwmakr1ktENU2nwm0m
30XiMVf6oAScCjqf8mp7gdHbItPi9AUjUguta3x0ic8CsAJenFVinnIDwLblYXCRyUSKDw+r4RiY
nIOVcMI4fx1P2r6Zcm/vLDzYxl6fKU5/7iCHXEHjBOrD1krAgZ2nIaqkUS42VHV9x7kY1bJxuEov
uAPYlWvo0ZU5mr5DCw1GISqyfjNQE+e0VOkbJyzEq+l/TKMFuHdhBhYtar0I5Ai7o85caw7nkOxa
oOqudZ6Tq4ynmE2nrJne5DQxLXqqmUYFtTwt7SzPwbKyiHRBs4PiVv5GVOm90+cjhAST+rT97ClI
G4mUnrNOiShfkuZjVTr0exCSD0rObd2TE710uQhuvbFXDN4hKYvFIoWQpbwvkMFimftPpXwTX9gp
/XXSpGWo9PlDFu8MkzTgstFG1uaZA1/kmWi6hGgjwWGSbf9959LUfrJzIuS/x2UmwQVzTDrZ0LUk
FUXJxXKe1Tq8HS5qat3SHmVQH54oLT3mMGPKi0riPXKGxleqNQj2t9zrP4ozbm6SvLfQOfC2z0Ei
Cx1cKrlDZD1N5slfD6SQaLe2YrpI8BraetH5zxaDKeOdoxOqcYE4Cbz8un49DUiv4mR+90MOc8pI
EHP+oi9DKNsyEla8DTMpuvRoSoLfRcHVBgDVs/RuP1fGg6A67pMQdViazWWSURyQ7x7ye2UJ1hMO
4LBIwkkpX6kvgVFTxbhgZ6w0be5hf/CQr18Nfb3roLgFo01/axUlESOka9kVtuAkFnA0iqNBXnUj
uf3HGYI6GhlM7PoMD8tCWa9X2weILFrlz5k/Kwc0v3ltiRZ3lFrykaud49PgtuzdjJ/K7qba9vTU
IOZoD1speCiAiEo+E2av1wHjWN2N7B28XZkTNh3BnepVZMivmnII6cA8AutaPRbjxuMdjz/6QTox
nApABINR25zshDKA7Hh3fR7OIfcB45lucaN8qofbOXAedvzWArCGsbHl3vpZs+fd3Ir4mJCB7OGh
L3NYEVQ573/hnpcgsKbfEI13s9d4FYuh2ycVQ/SxkT4xKllEU5AnZDMco0o5fjrJefWf4mZ+AdFe
/lxl83MFV2n0C5pXQm0hlKSBFnxYMQ61f5yBGE3fXJ11EzdU3HdrOxguJhe2KYF88QYsEol+Km5O
7tvVUZslls75wtYzNunPWdrV028oZUT+V8aCQSPJyj7oln5IFyyW+5I50z7Ia0+XN4kyKmFBkNS9
l5kmVkjFLRtOGOwEIIzT23oT8JP67aPuwNd5GkyHyBDV3JilTbs6eaJH2lcT2PuPYLtdVIx/Dpgp
95DZrArthS461QsBYFsilJw0ETCGWfccufyddaMw1+fXFURSSAeKcJAjPg7TmoTmLiVe9WtG/NIh
YVwL+7dYL8TPzrElJ6GRo0/A0B6q9VKP3obCeIup59ZzUkjJRk0a/ZILMU83i4uYCv5tBC7lYLNU
PIivc5xkEHA4MeKcWJMJMbVteJrOmrs18Yqgl+r/FDvX6tIfz94zQ+pmK1VD6nzKAX6mcwTMd22w
IN/H/UlYMsctORBWG+caGx3zJfDc7iWvi+GlPqGJWimei7jA+I7XWS0b9APjjKdbn1zXvyqPe/QE
yqa/Wx3hqJzWJ0dQK1TTrcY85mxxCTJWb49Gt8XBrm5BbXgcGjKvtYq2dUkUOhNZEcHeHdhqxkqE
x9kYTJ65yon4EL8EfBhJ+pBa7mM18sDW043tvFTvKo+uGA9fkXBWWT5WxaqfqwxQCRgrKtbbfY3i
ZO0+qxhHDVxS28ij534U4HWmJNY5YvaUF8NIdf7BcOHE6cJmU8mpMwp0tlPn1OQEpmrLF0xywqfG
NTZUvVM7+itWIerrYqXYkomaakd4AHGaRgdu8I0YRrPBL+mn6ksm1jetzcLi4goS6G0hppn45VuV
aVA/DIg6RnbmPh7Adm23zpQiz74D7OejUu+kisTPAvvZQNaVUfBhdzveLplV9a8r1ccEXCrp1K3x
R0HnmBhhoKPUNXR7UzWcMrpf13IwR/XOPSUE7Hzsjb2r5biOxy+BO3peXP5PBAHOoSVrLwa5ki9w
pBlxTVPVaCyFSGrHYN1NMNlLjAT4bRQ4qM+9aMmPXGPhTI08ln4+P2Gc02ZsAGN770zTF+j07T8R
57D5Sn9gQYvxNCwttZul3OivMO4CCWPZPL3pdPlmqDilMo7oEVCPW56OJrHJicE9LMBo4XQA+c3X
iSUUey63W38ccarxAvmWqJdFz+dI8z4ZzjGULkbxqs+jmyggQeJXNsA8aXoyDec22N0F5rSBCjtw
aHXA6x1BUTiRh0HXKdmZdvbjVNMzz9BCgy6EvgSSWMjbk/SKg/yVUglFZMytgT0SttTy/TxEHNoa
oY0oTh3CktpJN3/DqY1caekQnF9gLwIT71mYjiELKsfwecsG+PrZL2fS+h6WD2QcTlVHs57pLYcd
gVaA+d4RpiuM6W/+ZXdigtZTgKYLoJU76JPUEpE/4tZqp1INk0+y1kqqu/PF5e/IAGthnrTjgTHP
ux9rxOAP59W6iRqTvBkw88pZzlp+HvDd6sDQvwlvP2vqkKYm9c6DkZxeAJQSViaXqJLlcRHQdnQj
Q1GjsrxNkK8ZbL9A279AnQ/YYmJuy5JgmyDEUodQ037bN/eMbWBSZ27+Pzhnz2W+LLIIkXefbM6f
27By62iT43mOp+HeIaCdNmQltSBjilJtAmiSyOikp2IWyM2NxjJBGmLGsIWqIwCd3Yx/nk3CDGNK
7AvSLxBJZj5j6uQ9ITFm0n2vBRcsJuUyBV+fbjNgt3sKnK+TV0g5N2aN8Bqo7aU3fwAjeMLVJeNK
RpQhMpMfubVJnZ/H+DOiHuqBa3VH3o+lmaFXfI2lo+SNZE71Pw078IBpBf97IIrt+345E1Mc9eIR
y+7t3UgJb8FrwVB3tzJdSYfplCHo0kIg0gi2axI4IzmLxULn38jhXdiXaZ3hi/5pm93kDkPUer0I
HIzJ/matQELJs5vSC5c2/YSvwiVryM0b3eXmDa23HWvhYaWAcYWgbvwkwGS7KucgHqtf4wq6fwnD
uSN87u13WVYAiolnlfPeVpR81rOIuon260J7z+sE0km3dKCjl6laDQNdUu0rd4notaQ0Y+WcJVVD
/VmroNxHBpuffu+8TRAYaiSyvBVi2SywCdWE84C8LQDOnoq1UV9wFHvNfKmSkmsiXFWW69PN3ikt
1JJTJZKcMcgkPoNO3mf1HxhQYa/pC77sEI42xR0xqfC7fBRFJWt6O/dipOD3Yfs087IRx7kICG98
3QX2CtjfAr954hHpfVFtSc7ordrC4DrM6j8iYb8gH1185PpKBvVK5AGeiaCvWEkoZEqOgAIcpPGP
ojCNCMf8ATtVnJhI9pUu2IVDhi/cEegPV+wUz5+9l8NhzvnciaWk37T6d0u8n7RvydmhKe8lExoT
/UmcJIu3lhdyixFh6O+fiCbeUFLk+vXOXCK9/ea8fjfkPupgGym3tosbXWpmynE0xm6lJGGDtcHV
C2yTskloApvPMlmB9fdeokAlCNzKnwnNJZ76ZvZi7pUnd5oHtgRicJjpgG3TOiOQAgsPfRhjjATA
CxVBYooPyjqJ1D8j+XEQlXe+CyyvlvHrUMp9H+d5MesyttFODBFM4FK+4Oqir5tBc61DDGfkIvNH
jG0nXPcqPGjVBXuhA9Ra/8Fom0ChP8VZbZ7WDCNZ9Mm5RhoEUgs5p30ISIGVeIlItpGQriBD8bE0
7wprHESJzxo0rZZbh1gy5HWZQAJcevX2TLpsLhjCH8M2mP/qTdH8KwBDwzYGBDInhHth5onPRy06
n4b24KADCSM5SosebLEInndBURibpF3XYAj9InKflDie8EHkhT34TDVtxXAwRxbZqu1l2P3W82um
gjT4VbHDQNkhHUh9lD1rXrbaBn5/YA7BZrHd36jeZtVnv8jDX7QVpq43zJ+0T/4IbtcgIUAMlCxb
H1ziUQxp4JplqROFR8LYm2QhxqxpfwYMbD2swkm6oN6x/W5A+TqD57nKEAl12dEZg4mg6NAfG/zy
yofSa8SvqDCofA8l+kxkkpTILgOwA1c9fFtXKuxLGIPD5u/md5FcN6buG2PlBM+gIrfhbrsGdJhI
u9OAlQRxvAFmYCFJUQCkV/xSBcAa2Cas0zCesHZkYnUxHvAsf4UsTdXz1xVgGKN8VL7J36Jo+Tbm
hx0K8UPwfEfpH6jgYpVd5c10pfmdMYIrxjRYFePa8TVcEWK4sjXHBdjFY7FUg9ENsVzZSVxkTZH+
0Mwz46Taf7AwHveWPiWFHRAWSMT0MuP0ZLq8/X8KCjrh6+jd5faYtmrW737/lTmgyWxnj/4I3eyE
aCzKgGLbJtH6fOg7dHArOtnBdxkFsgLzP7MXIveFUjPmbbYCmwsZu7ekunvKZVe2z0gZ76kMxxUq
laIElKr31xRtA/6ZWGz8jcbAQfFo2HefAOb7Y/kj4QKzVP5x9oMd2CBpSFkbE1BKS6cogvb2pmbp
DinvaUullGR6+07ySu1N2a+0I35EYZwxmSVYFCPT+Sc/kskiqYgB9ZVbRf/mvUoT00jxXmzEGA4z
4fpj8fR6RADbUPFOXwncX2mzygwgauMG57g+tXggfEdxtRG56Le+RXt6nRoZRVKA3T+ZqgiAQHqH
a29n53psqib0uv23mRD0T65mm9pcZStnd6XqM7M4yhE+rWQJXy8YJ+SzJsz1jzHAws8hsmQ4QS4U
rvNgQ/I6AJ0Adg3XYxYFHlZL81WvbZtc2dj3x148IiKf+L7JMOiSMFDr0yWUnB8gTxCiVWCsbYCQ
xDP3/VyQjvz9W6W0vK1OtaLL2XXXJonUb4isSdTOXJUsHp5jcWSgnh0spKcwIhJfwC5hny9xqEk8
uLAJOYRU/q0nk8TnkrCxpYC6qYmCkAvkeTzn+HTCIz6W8/Kds2cadSGlHG1aN9Y8oJb+R8Fhtc23
Xt7xfkeCKWKtlJeKVjUypCzwimPjOMEMbpBPdzDQmJoy2oRDIX+NsX79tdmGDzOTbIAEWS3neH6U
0LbA1/92Z2x76G59X7kqR8Hp5ZrGBckPkmHXSWed+RduQ5bc5vbrWMag/3IRNKnsItAy7+v5segE
QZhId9V7bXJrae+PMDtbx0i0fWUxovB9ZP+w00gjE1tVajz2sUXl7rFZ07z+TxHCUK+yML1K1lWw
SePKapZ6KaMFN+8hZuBjuVb/u7+II2YrDhWzsYT+VjQ3rqZJ8M76qDFwvIumXh9Bbn6yjvKS/+go
9EuBbijVpYMpxYu+GXen32h1CKHIXrWrgmdpAvTkXwBcN80l4p3my5uLFka6T7G0+5yGiZYXrC6B
52HD8SC/HwkhyQc69CZo4eJzQz4xvL3mp/GnGrrFBzwexxO7TawW51DthKJborQVtCoEao1EY8TJ
eA16BybmLVYkSW/vNO0TjCJXojerub/P1mHaTxUxcw8DbypiLcO2fo/RjE1AkOsUzJHG7fOpB0qp
87OrsY23kmdWfJP2ScolrgrQ5A3026iLAFDe4yjsVldwKyC0UMY8yewSqHY4360+/EkUF5nQIXsm
9ju8nFM1FK80lXs6Ixk13l6ysUkaIWEHN38BKYyNq/2wwN/VgdCxoKpmRedfqgr/ZfDvdM7rpMqY
upj+aY08CSlB5ZnYHvxF/oemkHOYki6SB4XKWf3KbqGPaGTqND6+gUfkbWcPgDCcgkzSAcn4k5AX
MfAJ922SGy5AueNZ6YOi5D6kc+KL9w8DUs1fIZC5L2WHziixfkOl4oNy4N5oYv75wQk6yH0IdMhu
ojL6sBeqAgKgObX+VY5Gb942Mcs5ngY//QSMJcN2n9nRewEbT1Hv7b+YdT/MSSuM2gHzlpyZNfdC
VbOVZ003oRZ1ELynDdLd/7lRmWAADK4fCpK6+SbTi0bcOz2Fo5Iryy6ZRn2izTpVEXBJ/Xs4kTQ0
tvbgmPY/jxC1Yap0F4UlvUsurr3xlsC8yQYoF2Rxe6K+AdBIaqLTHoPeVYq3HSLzjROGTF35LF7I
2OHlSfd5H/sC53YJvJBpyythgYts5kvwUka5UbSF636Z2U5kVmlHntymE+kBMIlfd/6EpMSuKTP9
Q4g13LM17RH2abnmeyT4uzgoy//JZuC7tjU+6Jk1n62miCcN+KgDEa130OLZNIIBhZ57cFDqKX7a
0fBMr4E9BePNmal6uNmRPzXiUNAikmkwXJi8IPrPlGChTYQFaZkMquqGZJ+1wx7mSphC6p9BCHR3
ECuJhrsilhg4w3yjhqM/eNhak0nLU1UDnt7mOOKlydRFx++FyRddhR2bk2BoGxnbeLnlqDeZCIMu
5YRbqKFxjLQNkvgSY3k6qWABOCnj9liKvvVvL17jUTXGbSCO49/Mt2kuz8atboi3hyAGb7XHut25
+YgdHAfpcLm2+ty+TG1/irUnyvtkb+Q1JStpTMAFqFdFdMkn6uvXEGGk2rRmffF6mqOSVxiKfxPy
j9X5OSV86u25SDjS5k/ZnIyRfJX0ileNrA7tPmD010/7eg6t80xJdiUFBrwJRo9dZ2UgB910tD3m
uuS6M1SmT781jqjn1istLWn0+SkSYyzKz1eqvv2YAmRgGUrJ+8qsEAH6M/P8dLo5EF3c9KtRnXcx
ckD+QU6COPCZSRGoW3Po0+TYWhJ2sDLsDCC3YdB7Fy3MEuGu3PDo99XtZ78dH8KpRHDnpP7aBSiO
XoMhusnjPONip2rex5WoIKP6Lm4kAyM1XgPZeBf/C8cj4MQugMi5pQIZrMc/g5UjbBZQCwp4fjfr
gI4VfvCOPJc4gi7Vcyw0URE1TPHSI1G2p5Yu+bF5+XUP1+e0LLube1NbNdD26kqKULxUnS9xnelt
+9tvGxCLowzRriDFNZlwfTRxR/uYav1grUPpRkeJ2wB0QEa3ya3o/2zq/tZ3+FXCvO6BKZkiRuSd
CEPpQtQY0kGxrOZpvE90Yfo8uBK8n/9SYJX1r08OAOGiBTy8W37fJOFRUZ8xOkUxMtsyRg/8AcRw
0sOJUtRdLaSIMBoVLoQX61945zOIezx5dReSf5zA+6a4SMtLhoZQE5WjyQFOzXi/bJV1S5emjGnM
pVRSGRFHb3OTIfHd8nQLrB2Kj2iYfM6Bw3z1ZH74Rn7WskSjfztDNE+/HUkvYjZvw03yxGvkWT1/
16O9eRjFMKq+zou7kjoi2ZUyln3F4MJA2qeJmNyPKUuA3wwvjS9v+aCQ14eUZPErTbCbNiqqzhhg
rWF9Dk0Fguf8CK0bR7iOrPQPINg5KDH0SRHKGHIzQnLV50E6T4mDtXezJgc4ZjAabWdTTi7qT12m
6aj5S0WZVLCmVo4XyH4GPXGERyBQrtmOz5ZY1p5WGwuJHhr03LLJG3ejveaM7MoxGbB/sqIP5DN2
/+uFp7qS/YDWi98vaN5iz69HNa0V/fPqMCna+qNptwCgdzZAhu5n9qmxlNBqn2PQVSPdzzENVEy3
/IDS/1ImcsekOeBAcpQl/QrGvu0qamoBzpUF5d4W7hi2Knk4YT3vZRlpV+zyhWPf2YHxibethnfz
xcKceh+2G0gdIKKnKzewdiwJ+3p1Xh5Bo8x3QFcajmbWzDXxG2k21ZYz/q/kai8lsN3T9cgShmCV
sehjYR8XehdTId3zbcau5dzxpS+G0oEydiFs7MoWSR6GZvnuO3adFsMc15JYv6j2+uzbB+Wdx9hl
UUb0RSIRtpPnXH1DsSeSEloPNIpC2clLGi2wA7A4g/tgDYtOEqaSS1j8uLKdWkpfeIICkiTyDNIb
2xiy61nhtgYvWh2PaHZtI5RX03yYJ/fmgq8h8DBEJgy7+HaXauA00TgC0h+P5vc3l+OtyW34rPDM
BJ7BKYWykW38f5e1QAGt9hn2VW3e4qefn0oxssuPx8EPhSQoIz1lgJNz64u7TbP59yYXsgOtzONN
1kmRXkYNiSPd9eobqBhlvqneHP/UkEn0LL9NKRqZ5mmiMAP9THU2deihdLN7ZVslUXGmIVEN53bM
Ebvmn4SScCa5rtHwv5CIDiWfQ6QqRaoz6vPD6PaKtt1K5/FzrAsiOQi3mZVWqb+pJ3K0kNjQzG7w
NgbX1ZKcFlohmgOk890jeRA6DJkrcFebPoox0dOR3RbsJ/1A7PFOdnNTcPfG/xtn1jRD7ViWIDgb
lp7b4421NDn7OBwToKIceGA1MPtS3Zr5RqSDv6KKATiqRNH3eD+TKp1GDv7sfstOuzRWJjlZD44Y
0n0yZHmIptY0uZ2BQpzAOPgQuxOlg9wYyMU3aLsm9uwv2XPqvwd/eVQb/v1VTwxeM3LWaD13BSl1
7PCHcQCshVttucZ/awtj6XHA9tK8j6lpSEY6oVv2YJc7UKwGv1lL8IzVAWjsBJ2ryX02tKzu6ZiE
vmsEhIJrlSFRMfu4ZieEAXXiCDFmEzBQaL0n9VEHlRCvoxNq50HM7ut2rnyPIw8HZKpx8lko6YUY
gepYw3O+IeU9EUpjjmqy0HgIDMNxG7JudmEzG9XIM8Q5xWmp+ro3Wz7BSbEhY56C5Xw6zHiBkmlz
phCg9xNmJq7wIN+WCiMcPVxLSyKcegYfaL5qPWicHDwhb7uEOk9BlvU4Y+DSTcpsJBNJFEFknYwu
PJg7ZL0LjpEWcLc65C/2u2p4edlm++fw//DMMjxz5pfZ6DRQqJgZjdfMwHWRzbNtMhgqYRy15qnF
oQ75mkRFogjCVgbdfNUm1GlQ5H8l4PGn+eQemcPkTUcPPdfhfmn8cfSwjVPkywg9GWEeVRTEiRbk
C20O5fs56bODPLZ7F/R7ffgdosRFDIyunkUoVykiYsCZNf83JiX79m5hynwvgPFvG0vSjyq426+K
mILN7W00ojGS10f0n5F3Cv+DpybY0V6QPLzhQ4AS0p7+/NODEq5A/6xKfm2o+lraX3/HSANfC+KL
WKij3RCvpoTrdIWxaE/kA22OEl7sLClmuQixO+PHA7FhpWVSibeSejqqx4ylmCnP85k7oyiN93gS
KGWz/GseRK4UzNWN18B9mfMck59PCug8mFhG7eWglImVjeq/VU+mXMw1zHfpx8lS9/y5wk/UgZtm
ZmMSvr87sL3uNaPre1S2QapiHOQEmC9fjr+/a4k5K8RsZAHSAzs3fo1OMhR8d1JvPPy9OpHJK5w9
Lg11uURXt5uKVi3NPajX7FPximf76+hCoAzzRXxQUX00brF0InLxUmddTuUwfEbyW6t/N8pmB0LX
DzTTyvMsZfDW68DW5e1loIsN2RQ9TvIEZg/kMQ0c0sg+jRPaFbSf0TEvXGJmGP0FQxvl9lNrs/id
33/F0J7NqgapWyH/q1DsvmjigDJQn5pLz/8j6Pfg39RV5qZ+P/vggdNhi+Ekdmi/WQ7tJmOUeihs
rN+fSF0fRQpWpWQrWeN8jlCQEVXYMCWmXCf1QpuNnUC8FlFK7/tiMH8qeLGjCJ05Cn8bGVbbjk0g
CfFfQ5j+f5sU6Fzl66inkHBgoEfJQ6mDvfe2Ym1DIo0qxI8dpIJwZcl/Va+UzkHtBxlyvzQUIVwS
ACs3jnDnMrgGvH/+95eYSUd7CrafSiXN/du5j8+qoSn/Di60IsH0v5qYrRCfGmdJV6SbbTPQRUVn
MkoseXVyqsT9dVXmsdoP0Oyi8IqnMrbF3xNgrJvcPFLCZYXFmNnTjxw6OFaIJxlBDmAUH9eMQOtA
cD+m53eyHvJw9n7U7umuHYhJZFnyGhLbYgy+lVNd4UuxIwxyd2AUbsUDhvor57ofzaelyAa76UNw
N+PSBuVQ4sEjKHzhrKxV/+f2qdrub9ZGjwiyA9PtacpaZXQweG0vcO5IbohWsB+Au4RVvjThZS7q
4tMppKmB5I0sWVJRoQyR+MefkuwHbv9/VUqYvh2LoAmfnUMbyQx1XhNki0VT1NVYUqgjFYDH7Hi+
RZmq9ULD9FWd+ftJkfEKn62xUnUY1uM+2+H5yzmiOksrh6hS7JS081UfHSAgFHE1uI1gf9RTsN5o
/2Dtrg6MiyvGJv42ChbHNmDwg2m+lCfKZiUVB15H2NyPV9Y4DtyL/tITY8HQyF7ZER/5qbHIM21a
hHfzarMuxs7zSIFq20e53J+W+dAoshuvZaNnaKEGkR5jbBPyYG8Bhk91F44OvQxuio6n/hGwPAfZ
kTMrAb1qQQHGY1GB+cu5hdWI7CI0HmCRNpQpHMyG97YR+/Nt5Yk4ApB4ZagQ+psK9/0lr67Enpyl
kTbvPbwCLSrLN44pOxDOC9wZrxLnYmHVhFpToAQ0gvp1dgkk4oV8eDpE1+yriBX0CnKbMvhcoABP
+rPlamoJVFQj8t720iQKEw0vLZJaXuzFqHQOZy0nEuYObsJrl8e3EkdZyY6yrzwV2HyyCI+A+4Xc
9eqE29/gwwR2MXHFgWGW4F9wo2m2vSEznLn8boNOMj6yu7FawLikqGvz+8Gv01WAG2vTzd1wqGao
y50nByecybts0VYXgdlHNPuRn4NsfqDYKWNof1XN5irmcQi2AhnlZZi9m9J2/pX0FWTY+6ylOxs1
t9vfmfPLBAa9hU1/73ak2m7wRawg4RqknQ/h0P1kpg9N4iSyfj6CFzX/cjIAYsyI2IVqCmpC64FG
q7WwFgzgTpZ4C+uFeVOhdhXAQeR2jvm1BNvmLNIafH7R/duznX+IrzsLMOa1xKVPTWsnfK/0d7Ic
Ch4Q1iwCuiIUC50llT+7BwqZN4YWA3PraqpHavqphQ6NsuMb2RonL2lqMdU4bMbQ8FlksStxGdGS
xm2EiF3Yepu2I4kueeQ1vBPlQh0krogEpej1OkhQ7JUo4r2yrT09ZYxaHOo2Po7/0XV+boWuIDCe
1QXPFGOhHEcYHF7vYfPZsw4LjgI+nEPph7NrLkC+yJjkGIBZLbOLue0UJn2gEU8GxtLt8jwoU03d
bHIKjoJBSaWcaUkLUSmLtLbVo6yuTxEKzATkP0gAbF9TiiogZkEUlwRe7AYxXDYvWZkoAz4DNITd
MqYgHOE+gSvak0kvFPx5UM397GFfTcZQq4Us+V7vQAXEdB42RMDt+h51wdxwtonFSgwNsiSM+Q9A
3b2zPQtBr9YNI1NZvw3wyF4tRMHnGzmj2ao0YGs97LMtX8P97xB0TjnLQn9lRkjdHhtDR5WpafFX
ln1TqAtDiOUbFCfHU7VmETjL5HcPmh2NwuDNpob5KnslLj541R8MPqJHJZsQeNLjETFrmfRIGMnQ
fIMFQQLsIruk955INjr15RxmYrHI6rGJuJU+8y88DvTncn8I5k0NsLXZVOnhlGMlpf9GDpofpcNQ
qLYFoZcjt4oa363R/viNVgqeKLHRlW/lMZz3TR7IHhW0mtSvqSeGoYB1qc6kMBBsS6K0rzr/myUe
3qDmS1z+T7yuJ77tXo07Vl1+aUN3fP6ys+3nzOlGY/g+vA/pdKwX+9++osHeYhr8QSJxLkZAtinR
6kMZrX+/ysnX91EJk/W2Weu2e80mM5ef2+weu/3ThktDPmXdDT2dI/O0+1oLRxDWccRAABzKadEv
BgAbPOqbtep4gxWho5MQkYEPEA/8eE/93cmpS/Fb7p1wrGO+tLoTCvnOexNuzwpnGJv3wei+bqNW
coB1vx9Tle/Th68j6kJsmUY+aR1f6s8E1ZW6TdSKzI+i0hsIJv2asEPbIv4fvoXhmSdjQwci0HL5
TIeuZVF4FMjMxpNXBfmhwaznnOS2xw+FaFwsZNjEjl22ePGdQxFZDAtgeA3H+PljEtJC/LnhZLeV
YvphRsDMbnEOc7GjTBCA4FRt03Iu3A8beOtqosvyq08gdvp8ttp/7Zh7hpJBMxZ8MKmtqQuAqPb+
Ircm/G5YfFTnUpelN4M7fhkUEurwyFUfhGbBqAV08zc2M967kiHbZdmWJMVS+4ZVq3m7V0zaiIyf
WblpIZTwnuqTSorVaKp2+CASW6UXs7UFiW0Zohms5XMXCXgYOzPhGQ1KrxhBOmxWSlWFc9nxzOxg
MTs51u0dWCOGqU8kUU1h3LkQbcBOuCdpacKpaLPSN5g2zYXW5pIU/v4fMrAvXi+fVg2RAXfGRfcQ
/xTl4mNqSEelg1K3DaAOvTjLy7YQa7shVO0gYaWEi56GMXcdt2SlPukCa7LqF9GjlSY60D7TP+d0
Hzd0sAhDIq/5ZDBlHYTo+Haf5aPYqljzUXwuOUQotXYUOipYbBFHQYjpynxeWwUKlPhaDoWMkNpy
DzAQ5t/fyamWZdoUMqAxzHlSF03gPdYvGyqggJbWTdQPGVBr815sc0edhvKh+m+tp/iy7AxrIzZ0
VD1jyJDH8BKqK7HvHOvBub84EaONGjBQca5/xrRlzds0J/xBjdeJYUDJzp/w2x+sIFzGzjtyI3rx
+F96yeWMDbV9bvS38k2Uj0hs0icW+OawEdQVFxRnyrsl6xV0pWJoHuDbnzhVeBJPRIkLgbqYVm+H
/c6Ght9wKX8fHmzui8ngnhN9ivs+8TsnYDAN8QXGHZyudVPUvZ5QDAv45C495PEroGdLtSpcOghd
9Fov698IWm4ZTV92HFU/t+Lzn0j5bDONlDkHAplM4KpgwAmb0CT7AmbF6gclWLzf5G5rn/v/Nk4Y
pQBU8ADNgqbPtzs5OBAXLiBjv/N54l9d1Wu9TZg2LtLWRdT+6VAbi9Q4ti3E2XErPduYZCiEGQqi
AjZWbNpiCuWzRTdHiaHa2sRJWsbf8xvcNJKwCKN3MQW9gn5E4i4/fwwwESdUFwtmrWvJp2uQ6Uoh
sWPEhfG9WuB6kNoLr1Uc599zB50LVEww2vCC1u9MKJpnAIKDc3HAY69UHg0CBJg9S29WP7RE5c7R
6YhGgbdvVjlhwTxxPODZfaqceRCOyCBozhA3zn7yzqVhcHrQCq4Aq40l6kiosKvrYdmZrLCzxYNt
WtXFcsDkPtAxbrQNS7dp40LRCpz6SiG383vDyhDAdEHPriqMDYEp6jAUUxO+O4n6P6b8QDw+Rol2
qmf3jApW1ugVI481a1hhgbVrS9oMndsv05OAtIhyxBaaq+EB04cthgoPJmNEVJjE/vQYjaQwhxnW
3D+YsaMaBxO2y6e+C2fx+8KdaTGrpQ4ExQcGPPbbcrpBwLldpxzmN82tJAV4FiKVIqRnVETexrnJ
9Mi1gFENUmTkb2KC15rKbnj9Tr+r7zpFmYsVNnlttlvuOB1bEuYPeeoiL6zf0h47WTpc3Ztm2BSN
fMsDVyq1Cvy4oAemReYjnbjyS+7mf+PDNKQq2g855cttu2zcUKJQkOPh9zGtbwJ1MVYzfS6LvefL
JtJ9j09L4A49v5XFx/CNrpXXvHisCkaoIXHai0PJGOKILklXMZZ7uvV+moKTjN0ZQCJvEsX485H7
0YpWfPH8eVsVqgTCOySddNhDArbvgRwoVT5A84ArZ9lIJEDf/yd+KGpPoxzZ9bZMT2ZuTpUW9J6D
aWyGjxKG+d9HqFf1p3d1coEAlzP5wABtw5Jj5vU8CnA+X/V+LzU5eNfafsFDCLI4zmvw4/6nFMZs
ZH0rlJCSUQSLoIdsjAIpFkVhLbWxSvhYQgynZZmJBW31v518Dc4Gnm6wa4mk3kY5v1DXxC/N6gHG
UGbDzGQV5b054tR2T+0iJLwUolNlgBJ+YdsJIsr+pWXWpmfbaBZy9rlbUbK5hcmHhIOTT6zkhCvb
1RlAo8mwXYbhNV3hdlzXEePnCYOdXMR+8vzhbp2MfZSatwh3dld7ej3T/r0CZG4rVPLwsQch3wpl
Qcpj6ZcO8p9xJ9FWqgHGly3VbNLB8tixgYHb2ghV/qm0NyVTK1qztDpLASSiCKN0Dvs8IxllH8MG
HIW2569dQliPs9EQSQrKSEf1WHRjbTt7s43DyQBcQaLF6MFQof8CYj6T6RAX1jFv2MHpAezRsRkR
G0ipNf4QgPvCMAuehj5rgV1UgT7r2q7k6Yn9y4BjchB47acOD7ATv48EUIr4svb5jFM1UiG7zqUg
we+emT6lsv27SANrFwmF0frOKaytwKWHRa8gt/NgTQHxCS9l290r9h8afs9JkNzg9dnfovdWaMLq
iSxhgI7pnT6uPfUn4CnibvJQfhlhAvmT0AwGTaOn5x6GE/5ua8kxqN+gWmd+hmdL7FcdaXRglUSo
HE3u3mrVzkmtXGYLi141a0NM+mH2/80L5E0RHZVQWWKu91wgJhUpnrHDUUW5DKvEZ+RV/lUE7z2L
In5PwybD6P5epkC6r2go/26AENXlSTvO6oq5FhiQmd7K12tJHEVY8rY9w2EWdNui5+tMXA8zF2Q9
/boXYoSWEv4stg9NDNbwLIaTpHSQZVq/SERJ56ejqGP3AV4zDbU3Rrt6vWlT0N//H5+wqibpGSk4
2HOm8zk5fVX1O0CsQZWQpetQfVbJ0WqH1+88lGmEZ4VFH3N04amxJczeWIk8lpT2iFFDlPwfZYy+
fZL/H1VGipMFuZMOoSD75ZP+GV6X30g9uTxnmwYZp8KPMb5mMH3dMApz8Im8DqBG+Acr9dI40O4o
Q46jaHxlF0pfJ16BoRdDK6NFsAq/5rZ+kPlPl6LOfLfvFEBvXhKwt0Fnw8wllyooh+zAERWfeYkN
SV+dbvVBUA42/cLrxpHjpvl9aSrI3/W3Cx9eu03igzVsbZpVFhXLNuk+8RvXlnHBAfz1/db3xEWi
75I18NE0YdSzLcL7b/8lP81Hj7X+Mq7G2s2Bllb1OLIGH2qJL0TNHHkb+EXqR1p3/zFW8+q1B2AL
vYN2kis8whM7VuErD34AovdsLJG5Yw5RF6TU7+QVwXVBdKbY5v3t7cRxehdLk5/8DhqCJrJFpbD/
f7nwQdAyjVI35h/eTFl0fo4D67p8RGkbBio8gVDM0RvKind311315ikdKRuVqHi7XQVNVtZCNyw1
vzOffXCALIUTOrD1mXQx148Pt6PxLXdEqDx2s0sJS+6glq63ulQ8TRaZAvzSNjB9wmFIbV9a/UjE
SfwMJtQZOQJRc4b68FGyT2GrqRewHhFrPghClDv4x/an/rHJ0MePTcyoXzc4Pi0z8YMsW1aRTDQH
ixE52zxvC6no7GhBcyumQaGmadCXNLdOb2+oMI1+IUxHaBigCAeDCPcVzoFKUxkjZuYkzcSNycBG
WT7yWoCS3kUMTu1nMAQo46chzxufWXoK6HKLZFVh8AHQ7Ltfhqn42GiMtZfT2FFOWlpH/qbuXT86
SNg8d12UzKaBXF4mwvVfq//+AFcnuiGjlGmPiTz9V8p/jGPAj1ALiUvj6NstOFYL4Q0ToqmBwAfM
A6xFs+XyGSPUvbQZXsrgMPrGZOSdtqoe9Njw4+2QYU9EAmCcgccLU+mU0A2+vCk7OYWmkqlmm/VV
eVFBwaorR11A2QeiLXbMFEviioAApq2AAy83NHgbtMX5vbrYyLTCZEWab5NM4TqDYVwRi+aQU9zm
4M9BUFLHjCZqGk3ZRebbjgr+fCe73kHWFL+mdEaVEjQHXoMDxtlJvV/nYxnFejrtw+8OaHtnvfoM
2yuFCWwNcY8h/J3dU44nBFRl+YPHaKwlbwu6SirAQ3NS22ZezcyQNA5pIof0ObTotNSSafmdlJMw
lPh6imCa2gp6kc1y80PfeCafvQ0AmL9avasLij7GdCWMjs08Qexf+YuItRvoVRh94tUJ9ECYQrgV
Qj52Y8vE2pbEtAujmJ7IWq1LokEmxMeZQmjLR2DuE6V4aTZdeuNGGemOc4AVLM6AvoFMt5ScBYB9
0a6hoSuaLKq/g3tCjpQse+U+cJsrMDcpSVNejq2PL00OaSIu0UYnfa3D3482WaY3xumwRmFWQxOM
wapuYd58BmolJfwdDzGRxb7GuWOA8O+JLxDIAaMc9GLWWpPnhSi260k2te+ALV8ol2uw8AlIWjDc
su8LIagrkunHQSqJTlBuLL/wBZxZ4Mkxd23K3f707n8HxM/SqDDKOsHULtdQrzfxiAVo/RJklR2W
02M47HzlBmyMKkiURJTRBpH9DMFFkJicXiL1LBcWg13GXMoZrPbIV6jELbswpmbroVPtej+0t2rb
RDlpS4vT8bc5lzqyB/qrI6l+nenbTp7JgkSVTcRG0SB8g8lc8ctioScjUN4s0iar4x1Epic0qEuN
ok1qV3qWbAERiv8c51mHQuzqbBrBfkxCRnZaUVN4UGx7HmLPKf9mAgWNTgEoKx38htR2OSXnc4Y+
HEMuAg+AwADy4oXkqHcs39ky0JJ/ZZc6qqqwGZ7bhpWzDZgu5fn+p4fZNjPq5Yum6/+fbRIQ9GPY
bgroPyQXLLtcI7Ggp8tiJ181nOwESPq7LKa4Lm8DZ7zMBHgJaBcjBrxsi0+xj9LxUZ5IMC94mD1g
COu1Kj2DN5yjxfvrp04avNziwXkNcrs3iID+Nls56WmNQo5nlrTKxMmRY6GXM5wPR6qBjJxNT+NL
0e01a3NdJYJ1XzMfskL00lpn9CxSMdas4XdoAFW6VhDFWM8h9OIna+P+u0zzkXvDtFxBL85NDsvR
R6q/N7fjnm7KSQf5gt9CdFqMqauTTj1dYtsQ6HJ1/uBJvLV+ZsglXT5ygvFtR1npWQwBkSzq5u8Z
jzdUIqEeWyy+q9770JVaDAjLSs81HNespCe8oflP5atZLuvsF2EYx1BClg4CHjGyXiLG5+E/bzlb
bJC6IAjRyE4YfDOkiGJhgJHSUOuGPede+8A7ntxH3UA2N1ACukZKc6GLvE2Ajix2KbCc+TwFC1KH
LihWsoOio3DNURm3Y/kVPMkZOgN3D6ORIsUqMLB07I2TEXM/r/FKm0qs5jiPRuM8Em8rynmrVct9
cghn1V1bRL6IkA8QJ1yACk119ejz0ujLFujO1OAYVV+tyyekEQfijI4O5JMTbGTrRJ72i//eZoYs
M/fXSRT022WU54Dhr8XVuxnKeIBFnhiV6swABiqTejk/IVgqiC67BOUrbI/6dZZ7Do32G3udBC05
BTjksE4o5I9OJyK/xIABtt6fSEsinL89savVSI9DEtX7FPc6owiqzORhRbH/WfPGYPOC3dh8E+Ii
2aOqbcbnuzqSaQjG+P5KtIHB+gjup2DNVVLQp5MvCJsWMjNZ1jkgPfSD8ohE/Wbn21dafImq7+1M
TZOyG1qcmFpuEKUaxJTPG8bByiBxthxmp0IJeDYJL7DS6xmKvn97fLXWBlyjrX7KUTWUeSPHn4uq
kPAqm1sYvgbpwKNRxvdT2BYteZWUa1XCfcL5sCf/loGF/cpE285kdOZH/U/Wm4KB3IXuQeTWst6M
XSxBLmylc3FvAcCO+hYly460k8jiI2WlQLethvVA+0YxKUfEfyLGUjwSPlQ7oORTuOfuPIH/4mK2
7vnJWMAoLiJyATANReLlmEqK/8+kyvCDAqr/fQq3CzstVWtGPbSEGHJa2HDQSwTbE5/QzyxjaolM
5r3JWFlxANDiVZ1oB4JV76pwoMvHUuBTn9RKxQ77rnfWUQSV4XIJAl+hDBIF4n9hz8XgW+WW0mc2
q3EhboDQPLyjE6ZzAqp2DW9zUYWxvMD/hadjqvNInE/upyWiPN2SLgBnAczHH85fB0KSvdjnUddw
fbHePtaEjvDSKquol6uq6UwCS4wPQxrNJkMl6pLTlN2Rg0etu43ckb3xOkGu5rOedrDrRehkdVYR
B6eLvOeZ4VvWND2Y/LhyG3hHJVqgSNp9kQ7y23vEyWZ4eDeJ3ciUMHUgntKJRMm9giz+/8zgNk2F
PCmd967MpDM1g/I+FyhQrfCKdnRsswSuFZDC8AkBkQ/UmrDrwL1w6YBHT4D0CzAA+Kc+sK7kcN1l
8SiK9BZzY4dIfsAAT4QIo40r8Fsz+TFdKn+LIH5FUN2vtRR2O2BNACB8FZ3FR43jB7K9lZBQCuyg
Yg8jAt5o90QDiI7yt4VJyvjxmAlIZKqlTtyHoNWuRKOhJ0SBIzXvcHxoMPmdX9wyjYjXhfN3mLnn
wPCzXctX0N9QxBuJeSu8bgOxaE0l1fqXk/cSWReYL8RtF+x36K4GL1s5WodKWdMyaEW3pwFmOk86
8Cl5pfqx9PuQzulqWpu+H8pFZbltlNmBZyvSeTFFVpIEitIxu/VEL1alieKtShA1VPK3hU2HcfC1
XlQjFaqmG1E4G1akb2qKAo7l695TyT4RpSzoOd//6RCxI/KhoLYAc4RDGX3beEXG3dCtdtRIUomR
1PlXblN33ZuAgFAJrZmvQ/H3V3vX8atPC87LLLRP764rAzWHp4Q7JYjDayxdf3PvJlFGBUXRXD1g
KdFrpD/7eXchZNEVQQsaKNGjpYLkDTXuuum4XGPpTDoPJAcvkxwBBeND311lGszvQyETSAI+AntX
wFJW0gOlKX7GVcZE1/c+Qrgmjg4mzjjIHeHrtNUd71Fvqn3FH9WUPLEkegVKt9/n5k5JpiDk/BNV
cw4aA1+k5eegTUs9TQSJqcU616UbvoPHYYUwLUDS5UBpGH9D74sFzuPfMSzb2BMxytieja7lmehE
ALGhH9yHB0bUnSD0/1bsE46ESg04iHlg22PbB8qaIGPwWfMKQeVb36Z9hCFWp5ad6seUAVFNMgdt
Fcj3HsS8ejWbQIdbe6kZdEyPiUnx/RfGjseZhyg90hXvekC09PnCszavtIN7hboMjXEFGpKND+oR
xJrj46vq+MotLQ3/CG0J5ze+PLn3GtGhUlAMt90y3rG84pyZxTB5qLKB049CS8z/jBx0HCcdTQlq
71iMOCljOTJWwDkejG2ESQYLFS2NA3Xowtf1cf8uAsw4i1gC3K9gwbzS4cu5qi4/JE0Pu4j33w3b
sgSXRQ408DDxvEXXGLfj1FHSagV5HpF0binZRv44qzJMC2k2bg77tFVq9Nm1laRUGfXSGHQT3Tkp
Hio/vhoMuFATiMe6kw++s7AY1ZV3MNEjtSDSEc+iA6FjIip7IX6TVySUElC7Yr7hYZh5KuP82pOQ
YV4CCHh7xyPO/VMhjfvvKOQfL0bj8SC5uSpGUZM8f1zWtjXaiR30m8O7BmMJyDzCdZH97Cb2nsBD
DOdhjWFbnTU6LFdEWJw9TbcTPPtIZk5yS/17FofunAG8Feb0Okk4nTvic+3LsujD0xgtE4Ci9V3j
Ngwr/Ue2dqMNRP1/lGd3PCxI8IVQQw2rOZVuRKHuoF6oNSe3xf+Le8X7op55vGnIXz3crhaTNALX
50rf58NOjHAySZG14Af0HniIKHe2FIR28m4/5QJGQoW3PvZ6dmFxTIUh10xRAn8zfew5w2u+9Qsx
JEBliM0nYA44rnKOmOrDeURWiP8UlbqiCw35+9s4D1359RrlvGp1/w8McNxTI1RCP3I9hA70DFW/
XnpR3enZRC3n13IGuF1mzb0Pep+vY8U1EZsLjSpWUgstcNzhSEDwziLEGl93P5TfDk7q62P4obQx
IIqs6F1SJSG01ImCzFOsZtHJtsPCfnXmy3Tva/LqqrXob6supYqLNhKR0VwaO1a3drD5SZwDHpDp
t5baQg3fZIXeeutJ61/pQDEL6xODZDHy9UMdlFeCmrLWWDVqdF/pAvFlWT44q21ZPz0WlUGfr9k7
mpsxNYRTc4SypEOiHLUXJIvBn6IuVLoQnMu1eZ/SngeowV+JFnxeI2iKXeha+ALO3Y1AI0wNIvZX
QTANc9fM0E96Kb6wdvlvFBi7trLLyIABg3C+q+AyeTXC+eXB4qdK0G7JaB/awNZH24lhHvLg+1jh
j8+EA9XPzUS9oHeMZ2QFU9s+8YGKTgdseUr40l7kZlaDyd4RMdUPWz57eS/EFUtuBHTRnd8uja2B
nJvXlLkBGEKioOktQ13gGq8bI+mmXpQ0UvmYx4dpZSB+vc3UkZ8NVT++AMAJeCxgpLzFNj1tBl13
JLFfChepSXySNMXubaeooo+p4z6qFBPK/jrvvhiWK91vlVM4TpsHgut9dqNJDb/E1Xg6CIJodc1h
vDHv0FWuP9SijgihdIWDSGaRmXtNnpPuFPJ3Edd3Mi/acApHBDxqenXenAuv4oSrlM47iRKXuzlo
cvzyHYrRWFxW88RH63xg8sOnPr2X/B/hspHz/vEPr5UJSvGCxLb0WLBe/HI++l+GzSgU9WKOSpXx
1PevpmLcBYvKber3u5GNzHiTzaIlI17LKz/Mci+Op57uxgsCawNHCVvcRRPDYGZu1/l6l08rDk0q
93F2QtpBoa1F7sROxqCKb1m1lb7IqYs1jJrI1RQT8/poUW3bngCJYex978bG437w9CiR+zZxDj9d
pM/b8tPgKWM8SN3mUjjzeHWQwI8xJALhp6cX9K3Lzy7eXmByqophNRKoLHEkC02O4j6GzABwHEVn
llaWcnwG/6zNw9hoMdKXDeBS2z59OgJWSKbcbHvosBgeDji9L4iWy+sDuP5r/yK3hyp7k9h8H76f
Dos9nFuvzS7uQyPyeBS//78yfsg6t7IR0LKtN4naNwht5kfBHDOuIMsewMLcNbi0Jut4IiLdHgma
vH3KBKSy3oib2FYRQ/JPxakPI7mQ6fOB06ywg00hkcv6QLuD1w9wVq+uekhpORik+/fulGO5abZx
qbrHi+Qudi4b2HRjChVm4i6KAZvEio0w6WjqQjUyWS2p3mmnMuwvwydAvUfDsjuhssxx3tXYjEqb
FdxzxwIpxC8KW+YXjemkHeYqfj/pV9wb/VqiyT9LELyk8M6/wAkqFHF57NDYEL1XJevGAK0nbHCY
OaJqNiGWiDukp9hZO2qqjR5nG85CYAInCRrEm0Cwwu+JRlri5fgK3R3ePVnwhk0P3EGgGRwrn514
1dFvZMQZn+okpHUo+XIUPNWMRC93qaWIjnDbvmwdxYygVXim8NXDd70m+AKGOtg/SrjR6GKQY9v3
RYLPmoIO29j/UT2ZlZEQjAg3sdHqQBs73qDpjII2KYs0pXMgcR0ELrPn406ADPsFnSiHNejfmAUd
PQrFQVPwkMDIi/+KEsTs7Zjmupf/F+9kVt9HsGhRRTkLeJWNEWAB86kE+CQgPeD54aGS4b43CvF/
WLP/cIavjMzYzwIJpZ+gCTOI1j9K679EgmP7rqFU1Htj2NY13qe2YILrkDj4CRkyDs6cs7SFZax/
6XAcESGBKP2GiPhEVS7dUJnq4Oxj6uX6cVkoxLTUtLbzQKRR7+Fj864GIkBn9Fuzu+tQncCx5ehX
KCIxZlN9Gv2tG2ka1p74y7dJpNW1943gKdmbnhc9rpnbMxFdIlUkJJEb7otEOtk/h9A4i+RbiY2I
bcrlQw98GuLDzNutEDc4TVpXrC+n/BeB5kg1UxIXp/iuT0/KnFFIAyjeWtbiv0kNnsvHz2BmFg6o
eYaC67iSD2jQJpG2o0hnjV42x/1dF0h7sUOIADzGm9zWcgvY2kq5weyMRGQk5NYcsViJGBwiZO2L
/1pkCQDTcokXob/A34TB4xRw9r+oxS46vgaHhXpBLKIGBExZH4+iZOeAC7cSa7ZqPQ2fEWA3HyQZ
t0F/h1iolyMQGkZ5rxdZrzLK3zn/8zZUDWuYR7UK4xNOf7dL9X7XcQqEhPypa+EQFcwEfVAo+8cL
klbh+dByLAmA9jUc42MMMH1Wbp8NZBhUjwVDz1xGPlaLT2O5wB03vqWt1kiSHzxTGQ9AJNSTH0dQ
YlA193m6d55QlgOz/mENPBGeUfOgMFmaR6+B3CNOU4+8ieXx2t2LmEKfLnE9A5X5wDCFCXhWFccF
7iAMBHEWXZvIG5iJxhD/6GZuAQMHF02d4rgV7+7buIqBStsTvrB/uURwgnq6SGRkyUOFHG6f/D41
xAlA3ls6KXjAgGcotdpFt1oWjD/XPBH4HXMAipYPXRJqDhBJYejFC3E/Qzc4F3WymjYH+5Rh0mUq
LsLzQma6ElfzBormtNds2/E/WcuWkGLSR6IYiGoaePorBVmcz8lzJVK1yCn7kPuJ/8rzoM2Nso/y
aLYmnNNB9fV7LPoRQNCgEIuKAz3gtT6ZuFlfXhteAjms8IhsfE4PeYbnnqTr9/DxUCu4+j05/EnE
mxXo8JlqgShX6PeOkY/01XK4RaJFz1awtSpmHw7xvdEqZLxQBw4Z6ra7BD4qad5On3MysuR95pnO
FwmgYqgZCcY93KnxuOMiCkFni8BZU6+uja8m1CemaiOLkBVO2OQoTygPBCDF6zRJYXz3Va7KpB6N
8z+UX3v4b6FAJVQcuVgb3GdoWY0ijBygRW856uBD76bj2/6yIXV6QcGTdfhC1+RXEgEusDrqtYiP
Yi4Gb5flnkriNHvckXKUtXzz98AiihtwhKhYV4XdyRGJ1bmHZigTFswsfMJU35wvnKRnz3Yhgn4h
jC4+1+JZ+kVCy+tU+cxoarIzaZXahY8MJ1nwC5gJCzc+lGWanQZ1E5OJlv9i/ibybRgzbaGQIouB
514qSlAj/lRZ6L8IfIZ8SJ40wpxvnFcUfB7q5BBN3O86OQjg0xsj+QFjIDIPL7Ffeo4TZaxgtGZX
mrNhG+vZKjFd0nOcmEol8oQYxHblFbcldkseGFydAYN0XR9fQs1SKhgO/QvcKaHyLtPhgLs4k7DO
CEmyLd2g0UCcnC7FvcO7nI3WCqJ0MrrOJ1JGS1xOcgu9EnDKqdB3bS5ilTPM20oTKamdCRB2MM04
86VTixDyS5/FIaqd8nyaxPX4Eiv6FGKbBiYcD4lE4eVWguikdJA1dz1QzZSnWmjHzW3jI/8Oi5JA
J0x6XAeRIT/FQBZqx6A91LyIAawheEbBgVmBCaOyO8U/OBQ9gFHwtcqzpeA0uY2PxeZTfnAkJW9J
SDyKNPMvFJ6G8Z+WM4kMgrCGSvq79MlfbKNHOLBF9Ai/azx0Bg2YA3hTZXZnwhTKGAhZ48eUu1vd
wlCG1ZqCNGBNRdDiLg0TW4OPVSuhIqtD/JQooWqaHTlQonoyo2Sb8x8O7tKs9SYw7+4dzBl+wiUt
AVNcCB0vUO5NlLOXckZY6V5Ddw6TcmRZB4BkEbkhnc1ywSve/+OkB+qIPCJ8YLJmjrs94JVqeNm5
6284f4EvXbYwri8vupov6b0Ol1b2pc5vu7a8w/cyVopR9vapEASZ0UMC1+HA3fLRyF1cR6uOI9k4
DVivachpqdKAv/7EEttotJDAFoa0xXns/HJqRQVJHAyDYTpckRkyBtU8YnvTLX1TE5o6xv8vpDO5
rTl1G0E/yrqkgtG7yfgzu4ud4856N7Wc+BZF/mbsoCQ4O3cY41+zay8zjm46DVzcx/+npYhuuZCK
Z2S5x8UWS1oYROYEWjnYzug2aFbs7nxVPsFlAL5qdljJPj59AzdmsQalIX583KU6aUy7ntF/LV86
CbJzJnXjjVhh/uk1i45Rkj6Xwuf5E8Neri0Ml5xkaZs+op8kU8y5Mqiehy0Yra+zUch9fetCsVqH
M8yc9QcuycohEG0Nlnyylm4brWjp+C/d5WJ0+ZQMWqZguUiVKMs2Lf4A+GpPp4yi8fU9G0Tv8QfX
HBGL2LkIHVB+0HlsjZCIHx74es9CZGfkLjmYqDma5JhGJ3/HgfrPaq6AdpEp4BBNkeimfp7C2p71
vfziqczJwW789/dHsWI+ZYQqwv1uoCQYTKrImKcLKI+ZMhbqSQRN4lWjNn99Z8dih89Xul4l5NHO
52sDwMvbDpImEbwkznzeGTM+XmexTWTLgr3K8kIsFyDVYEERI1oGHAoylrvhce0+FsiuRy4XG3t+
RIROiArU7B0BGKojpQ3Ni06t/4ODIisu4+dchNoIQK22JwdYJ+3eeZzL2vSQiC1T64Sx/TRYaDgP
hnafaJGudJjyvqMjg5b+TAhM3rxOij31imjUH9WcNJPt+eALimwoIXe3Awmje+ha7vLe7BIFcWPe
05gdw2ijd7mnfVYuiqNkx5wKtNt6S8e14BLY8LRxsRHPtSj3KJd2qW60zeyKpUhvw26g4/bi5Ipb
kdcrGN0qqdwOx65zbRPOFn/1IN7D5+DG63/+dcf4/HxnTIk8dHnmK5NwOwXVJIPt5o0fOkGX3kif
XaJy+7lvHcWqwrZSrFONcxFmmHiJJwNkw4AXnTSPj8Bl0wrgEqXMnaJqEKpaP8ZWGOVk6jSrs8JI
Z+6PlHNb1LgEiwBOJao/LvMljqo0sTcAd03ZPfdqyB0O20kE+whe6fD2H1/5aSccWEQR5C3NRtqD
YCitR48lnN1WZ6B5eHzhkcJRA2Pn3GK2Jz/uSr++CQNbtigm0gJpBnewWYVf4qLAEFq3Vfoix8UJ
4b7iqoKHsAhGQG4Z5sJfXIkTPXRlygwLDW5CS4ymdEoYJ19hrRARq/bCBfS7XLaoHXDY6GET5Lmm
tEbnDKXq6cSFGcvZNWBcNXgzhQuCHLiPtSjub2Jsk2KJcKBu0oe6zPynNiTNO2GrRwwnFHGx3lJP
cfQzU4148vV9965esBeamFnB56t17xQSQW62eS4rEiyu5FMAZ6OoLMoKT2AJcf+V41FVN7bHBWbv
AvGjjgiJh9F8beuB7y5TBSpvpWNAfA/TJiTW4p5FDVtc70RNJVksdUvRb10nqaURy/gg74DuVOBt
35no2RKx4uNcC5dUsIHr4tTr0TR9bN/uJNmOwpUee6irUzYiUgL7YT9nsij4gw3E9+trRQnvIFFS
/9GKICZRoBVLrTo+IUM+eyWqnCS2mycnDRz1VCG8KvB/OM350opJWK8TAsPd//V3kA+gSTbPNHSg
HZLIDhwogDtsQtrXlECYrijULjcFJblSE91fAjLM4WyeHewgJDqOEIROky4BO8vvZZHPpF6YOu/W
7oHy8J4vf8RlJHUsjQjMxNs7pDLFIwvjq2dyTGFtQeut4kkg35PmJym0Ifj7ydb3K553kES0oVEt
5cqx8eN2RQV8eM1pbVNl4FILp2WiNEq5JU95QUNPFY2QhTGuURR2eQ5/8qSPsOmmvCUsKaE73OIS
ef0rud+SefqL77JMuaUYS3wUbMtWsKxdhPJ6Yf8at4tX9XzFKGfRyliWgdY/AS7LmPLxg9t/dzs2
Yb8aGInj6S3vWC9faezLRbRUhnPq020XEI7fQD5tuxJy+LS0NVlChya90Tj6tJhI7JIwEC+Q0Ncd
BU69tXm1C0Aklfnjz5Z+FLc1rP9KPtB/GMSqh2x/qI5J2TZjNKEUyZE/R8ltFTqB/m4PGOxrynvY
DHgsT7A9lWlElq+uG7aENe90sXQHkMkv6LI9xxkFKrVSpJrp9Xuj08kmK6u3g9GKZlG8NxP8UWH+
9WBnmzd5aPjVdFeg2cHeq0olEgP898GmeaZEmsDDtALK6zx201N3/4H4EXiACrOp3mEKtQo8IXZK
f+05qHlwhQ1kfzHeEl/l4jUJDtMT54UnO1h1lUXh9S7M/1gDo47GxaNKRGCRXd0kFZFCANyOcrBn
Fq5nPZOLjpSKuewc3sWW8YABPwT0ddrE5kiPLkgweUo4TMA6XhWZgMqwIHV017F9aSY9rDqpXSJr
o1OGLLaL/EajnBJtPO8PWjwBG8O5Z4ABVivGbkR7UPGM9w4nDdDUDVrvyT7hP/khijsPP1Gjw/hq
D3wNUqdxlGFcWAtIT1VYEullHd2/gbTJ1GA95Bl0R9vrHbVtEhIHWTu/Tbxd922KDimGgiFowPqY
2Oo0X8DJvAWNqR3vMuZzxBGX1ZhMW8fStjPTzyEinr9J54nbEo/IXEP0S1/zlPshCAfPZ4hhp+aG
GeeR4RrS2QBu0O1MFYG358xWBmPVJEWJ8JB6YyGya9jui9XO/+u76c6tRw8s5yKnmdGXF8eBaasm
a3DmGizyMbhf2stHBlk3bZhlu/WBYQQIbUkrnMBJUHHXAGHUGzvKrpICClIll8jcylNgxq3yPjx1
zCiQmV6EeRt/Jjm6RxOvbGfWg31Uh0eF/ZmAGguhxNRFtkLgt7Y2zhC/0F38eU6nGEWNQjST5TYa
RY25AjqpgMW11exBiY/wV5SwuURLqHuvNxq6VGi/q9CfZTQATL+jvYBVTRRgiUgk+KtBG3hE5uiL
8ZSyPPkB38oCjVlW4qIJszUKPzG6cxShRJRDgAzC61uxQ5RTzpulmTh8g775Z0Q0C9fQ75MlHDEB
Kni/75ay7wLhtB3f0LYfiAhqCD3z414tZMVgpCOyLL5/NoTxOQYG6O5HUrrQO2KQYL3R0lidcV2c
Wkn2SvbHrdtWhJhddv4GaU/LyqPHgPOB3k/MiYEmETO5NgAvwYVeBxrHU+5rF83eSTNmjhoSN9tQ
Dazlowe6f6grf4svGY0W/F0DBTXYw2JZbnOlUYysNDoTUwuk0YvBlxtfW/uaMh2AyodpFNwFZjz0
c4kkasdMOMUO0ZcQqHHLhod7L+0xfENR/C1d9Erhp4VwQ9sIjufWYhSgm9ZuSSOtyy1kLN0UvvHA
5iyEmGcJI/FfjwZPZAzFoq98nuWfZJCNVEU/i0bYB5xteDhJuWrF9DrXjZNLYH9d+kNe9LdhoYmP
NXIbHKH7Cpvep65On0oWJIqDuJjU9L85Q7W342l8kcHvXRJcxVcqYzsUq5PohQQx4yCFUGmDLHcD
kz3Ynzr2v8GBElwWT3mVQMBYDmea7A+UQHCCx/Zxrn7ZfVl+nGzzUmN/9REF3wUDH0RQOqffMeCA
DmfjpYV3Qj6z7xjwb96i6fC1rak0hAAGapTSe90T3ldXCkvAASjjtaG7riW4vwcHh35fYlsACwZ+
tYaQsTfxfwqd+LTA2vxA5MKUutC4KfezHROfWPCJJf/lLfywkXYhLu4GD0YQG8FiQ3qN0Wdefo1K
aXziQ28+NFVQFu6JXUCpk3kC+LrAOqgS5NUNp+uGbvMcwHImnsTIQrFewwz1cM7NYLh3s7ukDtZ6
DykTxnxgzBcNUJNMrx9+TpjLZgP9ZfgDqA3JATflD19kcxkNXkTa35pdMwGfSGxFKutrl8PWSXBi
ieU8TvegegNpehgFHG9q8b54QDRjnIE4w0BDxn5Xr1gREApyC5jku6j6+pZVPwhLzFmSloaVtcod
bJrSW56sTsGqFYfp+c5kaq4T/B/Cgxd0adg+A+cBlfQeuA9f6ARDz0OSyWgTjRPvctEQZClZZACe
wjk3tSe49OiZ6IZFr0QjHlF0e70Z3vp3lhTFyfyQW0Ry/3JMfjzUVfK6kOMeWH/Gdwg5JBh0Lg+X
50k5FZx4J86aWRsQ2luzuLr11WnvDCtj+vaIzYWqqyH43tan0M4TzC5fgCBAzRvKwWN4hM2ii6hI
lLrP4hv9ZZDj1gXV7RP9E1zkyOkPLDmGHD7Gu3e632qZhb9pSPQ329PvO7p4v0Z8KZLJnYqoZLNg
zo3KQrbciEqKnd14MCUXIeD/qlx2czB3CX9RL0xBzuvzzliOKYm1bkOJ9B9fqmhFGAnYPdSldf+9
VbFAgBKHs681atMECCUI+Jx10vZuIYyt+0hReQwPZfLe5sJP+qWM37PFE+SGDhX29GvXCI6dqtKN
bTZQa3Z9d7eAxz21tOQKNMJNXZtYoyegpYhGvi9WR7gVtupIZJANpS5enS+F+4BH7q/YDyFW9DD7
OZKcv7dvtnBjq+qNAgg5ZiLsxGnofTbzy1yPCI95bnSXJxF2mHuULsS16SyxAMOM5m0Ue0xTOZFx
9Hi4PpAhopiLoX/l5QcekZ8bjM5aagPMSpak93WiK/U/gWFOZjRRPDt1e0wu6qCDg6Kpfg7YU18U
aCMRyXShBCg2Ym6fthAROKbzC2wNXcO2YNcORsEgIigan70MhZBrhJF4RFX39D3WXv8DX9YDfAaK
euNV/BLSFwyE/xgudLIMGVJu+D6ocuzx69CaGXCDC+KGZePLoeK3ze4pvPew0BvrPLs0fHjKoDKN
+0qkgMIX+u4SY9ok9Siz+LjzNxueGiahOx9X74zFnvJ0QSEBjKdu7YpnrobfOS3kzxSEe8kJiygu
NNGR4EKZLl0TI74fMq7I/YElwNlrx4nCD+3Lm3Buu0lVeO8/KchDhMkJL8MLZUDCEVVbSD8IG7SN
31yRofgaNrFl5VoFAksdZX0MsUM/S9OrbtCU5mgV8pPjWSHLMwnKeMxwi4YtDwAdLKYvwzsxKEj4
Jl/f2jnfLGobz8xZi+u47szW7ISFIzQ6nEDfqAdD0lROD4zVuTJW2EVVVRHlb70QBQ1IS6kvsZ+E
A37y6H5tfzFKSSrjbG3ZUP+DRAkPuB9SIOXtoQydtg2Gz96r78Tf2tTTHCZLgCwkww4TjzLIuEkV
NjavEtAjt4RX0vJjWKwa4itbrPNSoVIkwHVViyyewyZJGMsfp1JBTMREWFhW36RIGBzznfgomicN
UdS8l6Vr81ACZO8bwu7Ns4Y4k6RuE2fPxeOBCkC3F1V4YO+JTTInn13CV304hj+LE3+7MHj2QGDI
j3pDQvIg/3i9psn6xxWigBqTHlJ83zH/b29c/Ou7ToJfP+nttVaOMrQpnJ2vLbugmV9tracbXBg9
qOZDdVdqvPFnN2CRc+BfyYjZ0EoDtQYRX6GQZRuekp67WdhldMPNKCFfUWCxe+ebTMi603W3QK8x
v2SxFr0t72Lwbsy1mG84zdkGo5R+0rLKsChSH+oBZ3vNVKE8F55ExTUUJbq8LANKpOY8RDkB+h4V
SlRXM+nXvud2ceqi6pRaD0+JomK+uPQFu0QjlTq7jV0xva6rTUm2BywnD7+x/VOE7tvd6JnUhzHc
wVTxRj9cC1hOm2mGUIEp4zjQ8UVUn1AGomAXfv3/qEf9nqIS+pFjxRCPKoir4JbY4eg9AvkkRA1Q
hKwLB0gB/HQfdPUEh3fUhAAfXaZ7GoBXamKvbduK8em0z/+tzvqn57atvE5ISWxBq8/BciH5r7qQ
TlK2w9CEdyUNaUaxDVN+b1iA4FyHboqlyb11B966R2cP/lt8Gg2stmgnodLxLaEv1F2IkP7JWc/X
4/8luQSYvrZCCwvkM80drAmvh5il21JoV6Wo4tCPYT/gfJfYrU53UCvw/GuRWFmn78aO1nj4H3yG
16YYuuL7tVcoAonhXxLPzZKbqw7a3jrF5oTuDjeH/zyk1vm2BmkxfKDYWNDCnsnSXzEaF2kEnmld
IVo9sVSL58d+nv1eggLLQyrVaP3vT49/ANd+qMzaDZiRpGEWGCdgNOUd6KRBu9l5Ify5KNNc6fnG
HtyojPLpUWRli+it1my8zSZw/UeO65CZIRJmh2IP6eRHLNqIWTNY+CosZqmsnm5+YlsX+ynWjYMa
uoJEaDofq20I2BaexZ9U3fjAgCyN+sS0A2pkcveftS+DkIPgaM2FaHGS5n1927/oP3ilCmCGikeq
bSSjOl3Em9L09/EMQHBBnrkODDcm47ZS88yovY1TFEHwuj/r2+dbcqQwYr5gyY2fjRac7e8NDqb1
SDxyGqyf2g3oQuFVtfeznF/YNyks9j9/8hQMfrtbrtDie33gU+ZL5RCz1q0GDpKS29oiqlHfb23e
D09kU8NMfVa1YXc0B0KzFrkRSMNHMcyDURCBBHfLEo9y6IuuFSSV7sidqaJ9Op+iO2aDoeS3/kah
agrtZgaTBYw2fMDrWfCKiKbj9lnVjsMhruhvhN24cdX5CFJkpmSYs04ms7npNm0Vkt7I8KESuJb4
DY7MarmqVuz0MRtEmJgwoyhOsk+o9+Vl04387mIkn8sHB2gygVrjSiajaivXSr6T2/Z38eyPXf1n
P90AO+0pD7z5RPk6sPpS/F2wiK1onG9Knm/XIzNw0GzpEoT6LrfRawLVQXyk/g4hWfy6q9pk1XeJ
KB4uP9DTh09fvhVcVIiUrvScT4z3NN76kBqfdpoukYMJRUPynjR+JoFVQdtmwNvnTGdLEtwZpdCe
sAwxnxmUY9CcwybzFQDKvkzvqpfmHLjj02+NVXJAzdkwLnjA7+DnkGCQFkms1xc7oB2lX+fXL8mH
ICZPV0fTaLmhmEITenvXzznwDZHIJ37Xv2hzifXoRzDl3cBuV10LCaV1q0zlqG9RmB2UKyvVzn1o
a6F5JV/SNkfcbsISw6f1Mg8FD1NmO0OLMK3MQMguqst73wYc5oD8ZJLUg7K+ptocH8sC9j5YpAJy
TRBYe5/G+NGT0xR5dSLmDh3jOvDnd16RYMlBZ0usV/eoZRyx7hu/Dfqzll6dwxc31F5DbHQz6NJ0
G3lcl6Lvx6bB7ohCtM+eU464O61OaoAx2qj4le8i3nyWzxPfTll96jr/S2ela5rHBQI0dn/NQ8ip
zHcuURtwGys+n9/e2+38VQTT7eyoLxZdiv3BKQI2fTIghUiMMur8rGkEn5cuPwGUv0pdvEFgdxj6
ev6dYYCNHhPckhEMTi1MaayYLLF0J1bHclli1Ttvv/cuZFgKYxEwO0gJ7/UFAdpIabRNn1a18wv0
AwqJYOa68gsiRjHvixHZOG6/xCpNMDCQAFAagOM9q9enB3HEgN1zNSLzXQqNGpPaXTxKNnOCGLfV
OTfnsXXs+chWpuzN5SbROCklFe+NuCqXCW2wsGgZYk1g01OHzEkg9bXh06Ebsry5naAGAMDtxEGw
eUiBPct40THBcP6dfFx+cbeTjhX92ea2lUwK9AFOtxf8gjqj3Z8Yh9eC7KE9osZM7ihkQFFbGG/K
Jns7+lmxSNnETkdyvClblm905gVvULrLDoaAWNPkoUFoerFj35yJ2Wpd6x/j0olqdA4zDPMLKWTm
PCaffagSwSiAqDwPFUBTDhRHDNL0Z1b3a31Cachbpibq8s0ZvtV8lz0Xv61X+ANO0WrVLFkO9c9G
7q0RSY1AkrwVcK7+Dl74z+xz9A12alsyjJsCuBI22dxv+wDNUGX+fYXIHv5rFx9SKcOGnUYd40yx
9CrRP/hJDkB/ccT2G8ccIGvRjv5xJX5lLCXsGaxc5NNb3F4oaJsWFjOhvR7gG5/fWMu55NaQKHVI
DBWHxeTwoVxftv8HeGAnPcMMp/UuECrSbAEcSMwPK9ffR9UO07t1HazHJmeIKBvw+NMNPv2tosY2
2yZrlIQwf8Xt74nk7Nr9EjWCBXhFM9HA1QnWaWJfrYdumzLBFiS624JHWjDr5FVr0L7u54il1dko
DhgklZ4X+02BMdKnUfuwyCB0rW9gHofdIUyhgreS0QJ2k4uQHAvWBv/5b1mJ9bt1ykzsVhNsWwRq
dTFN1UbCBmk2dyuU92XQaRBSFPvrz1EyiKPq1uNU1HEejphsf9KeZYO1piQJIqMAYksK7E9qCUsV
4x5KBMFx5ggLFsiVcJQLZpDKgbWnUwb2PTDOIvgIZ4o0lXimWUZJETSFwl7/+o9nlsuIBQXTeHrC
mWKKX5wTEQJPGhqREJ5+rMQ5cYMhyJGoh9m94R3jxOXjvxBg//RIlIMcEUYH/C1aERkuWqIjzGVk
NWHTKCNvC6L6HKD5kHkEIdpmj3Ji1/PrkABeYq2ofshFEVwyBE9B4oLkrh2ZIvBUL828lmNGOegY
invXdyKdzla+atOcjsXSssGcnJTpEu/mqpn/RinazJdQRlvm5VfY6gcFAGe0aiwo/SkvlmJkE6vD
N7aGdmtf+pQcRPeTc73Vr5/M5BFzkJBEWglraBVZ/UKllJXDrPdB06JEO2/vxQYzJHOpfUzHbvAX
5Qp8cBxou+2gdN6tAOYDLRYdREfil0Lt9yJWkyn7c4y14y7YLEOcMAuzov1EZRloMIUxSLJMIV9D
9lWwUDGxy2/gL3crFqi5SaXkJP9xQV+vGsXD0N51zVITkwq2YW7NdHw+5INU4Qr1BcecSBF+jysV
EA9cRBmjZmJnw+U4rsmDS+6bi9a++OYJUWlwfx6vfOiMHSg29afYlOkCpy5P0EFVz+6OguUn4NVr
lXPFjllymLyPgZsAds+OQCvzh5aI7l7bHe+VJpXEeCc8B9EUFlKcULAGVVcOEsIXfd6rkh7BcC3K
p2DMWwocdKz52bLgJuL+W1Jl06bjK3d7oSO4K5osAsYcZfQx0ow8nLFmQRJfBgv42m2CXZPnmUu9
quuGbqtANE055kiWIyJ+OSM/i1lpY/qDxmS4SxFS+c1sP4xwpTu+W6CUTZda8GgVsuDDUPNdB/Bu
1RxbfyEkK1WHSM1GR5Zj2+5GVG/AtX0iYJ6jw7eB5SLI99IuB/21qVXYi5R70MDUC/yyrqkiWD27
gkvqb1/boIRuSmdsVjAWwrDlTlMxlxdRnBwAMw1QTOcj71ORDZCXn2tl9YLIHpD8uF+wJMyk123+
rk9CAC+WxUt4Jcn1Gv38FBR1FOykpLUAlIKVSR53hMlhYeIQMJYPhaGdm9J2x6br+zbPu8HZkU4K
WJG9d8ocEPXyD84nzIeanSHD62K4VmgN15nAjw4QsWB5dKgaeHq+HA9X2TF623MkEkXHpHMzrbFG
wsxrAetp8m1Qv0jZwHLunLguXPCgpWsJQeN810XtsZdavGKPQJUQQI+1CTvVjyz9EOc8MZl//gPO
1AakzLg0i8Y0zcKuZ2jt3Ec/W3Q1TnxIbGccpfXxHCWfdCzd3hOcgcIlTmvXhm1BUqrsV6Qu16hu
1RGl4QvLZl45Bc0IfmyCchOgrsiT9/qJ0UmWr5F83KxfbTN7ayjO+IrSdGU1VU3hUup/bQ1FLrse
Xl5HQ8lP2DhluXOE7u/rGsZiZQ10rVB2F2z1ghhVWJtLw6g5UWBgrFAns6v/xEUGvomUwVpRbEVQ
rIooZmFwW2lU47MzMF8Vtb4QqgfmNnfsEuckgJzZHZ5N/i3Dl8EXoPtAoWfrSPCIeCQrh6ReArwa
JlQdAB2nCmflZvUa92Up9rUfKlLGEcGW2UfitJeyf/9pbRNs5Lsn7rXx9cw/hjGzYdCLI+TGhFwl
/luWsRsKD0nndMDmCK7sKYgsbmcjUele0o1PDE+iQc3GLvHcWK0l4Mzu8ussB7W77W2Krc+uOc14
Ok5fbGMORKDoqDt5JKIHFReD79aSlgZotCe8mxNtFLlFsZLauZblbxd9OaPHUG3WK/ZOkaJGcSgv
B7vHBcV43sW97Gz29pBegI8DDyr2CzhogmB3Y1cY+6/Tqdr0f75gdZhds8OMZBOMGeydzjf2ZVgz
h3XOSFyWhinTcphm1TOr7snuwjzL4TQTi4sN50x+DugBT6tU/1eVN1iQVEaUpktLuonqFY9PH6Bf
1Y+f/GRzvKfuVPTMx5Ndzo0iLrUA/QslElfMwQigY1ByUPxGVksJrvaDCIZmpWLHa6q1Eme5PUNq
y5KALDYhyiHOjRzZyHW0Gt23ea3BTsfMFlhIO1qQxmth2Nu7DHLeSkRyDEGwKSIg7dyUHu0a/Wp4
OcmT2y4IvcPpI9VD0EvZGPSUyWISYWyhSM/oibrjkNxrj6nwN/b2kxlUOQt4mpMmrNHrHEsZGYFS
C+QGb06kCyzDQbIRfZOsqkMiPD4B3kPprKCl+lpwzqwGMtpfm7E7loGuPjaw3P8oNDbC6qWfU1at
n1Yhrw2vc2nr0aCjUbDTXUyNx2ziQlDu2Wq/dgVnQUsnwSIH80B3llGy4mno40xU4nsWXjeAg30S
9cAidEjBAfn2hZHfA5uOLiWTjvXbR61J0y0H2fmTq7eW4HwEdpqxUofr3/ky8E0aXI95Tu/QnUnE
+H/c3CMbZna+YVoWdFmgJZRc7ce9M9/I6TLFuTNzlhR1QWV4AJAm2mM17q5kBzlVRPw+31HJ6aXK
hfgBpePAVZ0UH7p/0y9BZNAX9yQoDeWR/m+yg+7+q+ZOMQ/TgBOI47et9Hs3U+O5iMBVvr2mCcDU
Id+63PPZHVhb1eOAm2PmewjsuY+rclbSnl1B04cDuDFGqQj0NDu83qJfHqk3Iq7R9f61lO1u2/4b
RnipLqln+fwEL3Lxfg4g+P9+uG+3gUPmMXHF+Wcy+UEwi+8U6b7Zu0laLH+0R1srsV6qQbjlVq4L
oCZa3N5K/oA5+BpcN9+QLL0KTRRgghXCCtDmuUxdwfhgmSdS66tJSek6DlRfswruwKhyLuWN5EtY
AVfwArkZrFrlJu99pAfJf7kqjt5rAlFUxB/+sZY8rvhULoVme0C6pBfHQWPsDW2xsiKV71t+GPiq
GkCVxPGxJovH89vKV+8gkMEYqk/MrqJwURqODmTxrGLgQMgvABkVmPiDjnanAlmOQsjH6gK7pjPF
AR0ysgS3feB+L9TPrrv6Y5BDkM18/mUB91VIWQ80mmVxfZ8D8LImdber8CQtgkLBKlt2etzjulEN
ZSc290CQQiqJa2q/0YQEELpxs2aCoIDnMxrUWT5UopfCkoG4QJAPFSfDLmi5Oz1kkYhcDzs6w3ss
Covilh9lxr7H4gm1pWuy2uCXVkiKUcSC4PPhvEwazWNl9rqvhl0466hWJ4e828u+iypTXzCNx4UH
fx3htvIZVCE248tmqJ0vEBbe4NLMtjjvmu5Fr4QtML2VJH9+BUH+CBZunjC1xyCmc1TAuMgF5iKz
eta0pw58RqBsAY2Y2zByaQy7+enecI4T2DCliz9LO3+1O3JncU1NRPVAsyciUW2dcc+NanYJeQ2G
RVXlrQf5Qnx2rE7ZphmQbpDYj7wX3y2NU7S8H7zJMxKDjDX4a/iN+Ol+3RYzA5uxsF9FFVg3NxjF
vDZNBAOxSFOenNYyDaj65LgY3M3MGDSQgM6/U1E6T0tTOtooexARtahNQ0dnZOH5hNfxHGBC0KWQ
y9vOZg+DyuVs6mS0kS8bXUmfV5P8enPeKPkTET9/guwR87q43M245wyxLoPZ9vUvIome0dQ9jnWG
x4T3s8yGe5nW5xumicUHunOXj/8ZViRPBqKpd/3+PxzbPXzgfrSwS4c9Bv1Hj88hy84tPk0CiVFD
mm97QD9qdt2DPblj3X8iFhFJPmfCttwZBYlZR1jv5oxvyWHjhyJS6o57PCN/2Kj1Sa8tEtZ4dV8Z
Mv8N/ZMwSrzzMgNPxhb9qayp7Err6nJgSPoA8rSjkjqyZKvwzGcQWT2AAlaiuRasWNhhsbCqetDK
fMBYvr2tL9zuYEVaZFn+mORVN2xtbL+NZRrR7IlRlxYFVVKVs3W+hrGcsvm0MSpU7UkEg8K1p03X
r/vcRtVXJXC5M4KCUZ0Dbq5unhb8GfwaqHUaIHwjZ+KuSYgsh8M/2luH4zfDjoWpzCuDSd16ZMp3
ab3burHWeK07yZ9SaTHCFdpc4JnJNFShOkSzla7r7oboFX+/QpbG69ZVYejhfmlpO98PueDI9W8u
GZWOBTr8olDOBPobx74ldvsjofgR55kHa7orra56qlFT3UPnv2j00/CfNa+b2tSr1+xAU9z0C9pC
cykDQgmIyNUEBArxFj3EZ6D6KeNFgdbEUIWGYifdJsZtG4Yb/Id1oypBNd/9sEYt3E/54LQ37+wk
OXALPICLDKmL9pVYyJPj5c48WzgFiJA10AfXC68LOJMLYRw6rjhRgfgA2TrmD17+vlpU1PlUII3z
tunfZa8EhaJvpO+GDKHshCUuizcGPIAEYiWdM00n3c/L7SgSzgJaqvstSZZABHQf64otH9RoFmKm
FpZwo+m8w21T8TGiZ0lEfrzIXN4o6bsm4SHfhXRffVrax5lJwvf23cR0KyW6I9w21nL2DiH8BsIu
ehznwUGrjMS4VLpU/tXMkwUOkYGjh59nNAovsBrBcB/GpHUBGzqPWTw+knAZQH576rYKmX3rpUH8
V9CiMvEfIC7zvIwIvCVonntd7qEbFHzlO3a7pcePsas7Ns4pIBwTHgiOF8sgIu3fezIkEHy28pk0
MH9C7LiAdpWascnkZs+PB+YulBTE0x6gp6f/QHrHtevpuk4Z0hfFqtMwrUWp7q/NMBrm2FWCUoKP
edPsVnfNNB2WYkihg8ZYJW41Cfblhb+B1WgJncEW6L26yxawdV2DzA+Z0GTCEI7KtguWTBWw8qoB
lPzu+vtQMYhKrz5hIqgaGOKKthWgFXAPrP5G4Q4eAPmz8JN/xvyKCNc30ll3DnqGXJ/n+/6FyWvr
cv/UrQVCxKYz9GUdsNT32UP6DNNmxpCRE7nl1Aq52j6TY65ZjSoNx5SmPLQmcnKvKdKwjArxyFNp
zh5EGhplo6iQLgIq2tvOoq76Ipp5ilTuiqkbzWgKG0vBgy3CZVybcwzl4I9YP6r52SJpkIImwoUS
BvjaTSVqGxWU37oGMzwRP0ZMX8LOImD0pxIEwhR27bcZA6TLrnitWthfw7AzbwZ/cIN/A4nk9A3G
pv7DFniitd5HwmEQddjRDw0jjU7UYnHecdT4kbOEigJRo9A3QoGz5UV+j8xFtiTrLdc5EWPQ6SMw
gBKc1mPYlOBnlPZHRVWqshgRTOYWbzNl9s5fsU7PDuMnZDIQ65vWqEShFC/cg/MAil7IMUCVEnkr
MQd1+sqA8lqVFiBfTRMnxrmTX8PrixG43IGftXREls1rLYFRIuDg0AcAhGQ0j61bjCrn+aHGo7Js
2BXt0EJj4KDaEF/YI5wYF8Czy2QscbIqr59MuuHE+RuPWWIyAmlGpLDWHcR3/vMRI4OyAPIW5rRI
i46y3yteK7lXNUcl++Dl7OF3njQYVzxt0US/TCySRGofkYSxRR/70ItBsJ/R4giKyNPwF3Dli9C/
yI0Kp/rgcA0K7kHgjBwMiFmp4iBh22YFlb8VWegm5cF/nlVixjIq8XGHBfartJHtkbvH0ipRr7YN
NPtk/38gPNCrPQEFz/GNcNX+6ICN5eGbAHEFVUwmYwy8mOSJGa2h65ykLLnNiVGPKlBnXsZ3/Ff1
ErXGXw2I9ssDGawcYqQO181a8gGqfTfzfOkqT8pxeP5T3mZ2GIwi+ffJ+T0vcXPJ2LzEeywLcoL8
xYkbAROGdXT7785yXU3GH2ErZ73OFA9Z1O0BU2DsQVxnCv7wqhjtC3Ie8DyUkMZYaJczOuUtG1qM
6m+omTTqZ8h1KpN3z2apTouHiPbrhHGLjPCzuqmjoErddlRKtPoKZBUsaGp1PVkBKjjagU7WgH98
1FbQ4LP/hJyPp/l1yfDT533Cr4GdQ07yCwbUYgxZ3K/3fVsl+sSggFB72l9jWDsHx7r8JQANdAFX
iyzX5PDXY6/suJODuF9OOjEeczsLRixzw9X4f8g5J09LoJJMDyGy69IleuLZ0l01ZZNKCB2dWMIN
NO38OfPGGqZEvRg1PYZHf2av5UGccy2LSOAUNhtmdfZyCOqkprXtwC7E0mkJvEM4u3sjOj4m7Ygc
sRf9EKxXDYFQRL/9e1ohURG1PhLslHXEaQHphPNGnKg7yQm4Zgn9yzrSwPoVb7WGuOX0LyVa/iI+
3SWu7K5GusSv+yqx47NH8Rh/HpZRsYMK6ZL5ufwMezPfQlnErautZWUrppkyXkQq5+UNXdMoaeuT
t8vlHpgiGwM3r0EEeMXXDyP1R8UhXIWuDI/0xMpVam1e2v7zm0fbds2McltOQezhlzvc2wsbw8Hl
w2gz13KSpFnnrtyBQxtqLyGJ+ecEK04RDzVmbFql09GUlb2vlCLyf3qrOzoCxJUeBU15xKzAQnzj
fFxFePSJeGAFBik0wKTm16SNeozPnvaRTSQLORi9mC6yVGZCWZDfXwtYzksFK1DNmRSj4fNrX9cz
tY4P9FV2bo1ZMpLrNhokfBVh44YdV2u39CPYmdmxGfqPB24pxfjc3MbDVd3J4BP0/XxR429XEcwh
CJaZ9a2B/qVu0EbhEDpr2Xvut9a1jL2klwLW3jOFRu8giQRnoaX5F5TBj2v199qWW9MFgRXlIgem
XdBmpM+3oMDJkRYvAQ+7j5EtSsl+CmDSKZIDErlIcLoe6eS80TYK4rIwDIuZaoPGWN+QuFERmlm8
RWHhCKCHasTm1cGh9Ql6bv+pG9W845+Y4djZ5Ob8G+dHyVTU0K3TPmXC4pNu5dL83JWyacky35PJ
rGfvHW0VeL6espFIuiu8oV1fpY1/ZIMkgSDV77Ld/riQHFvB5ZOtcahlRWfvW1IsYOliIB/Sb9eG
8y9NNwgf9ZZyy4HzY5j+EKLFb2j1TQDYKxwxHNavxTzrrC4f0yTpnpPIDURjcJ1nOqV7/C1ItbhZ
jvwT398qc/DITCjU+a7zeXbDWGGUCISmdjNHM4v0AIjbDCKj6FcZY1GEUs4PR0FoNg/yPOgfE0IL
N57kiJlQjgpdnMBHyfluTc3kcro22HuOrsqEky809S7ZXCoAqZW6EZi6w95rOUfmdlNJwktAaf/Y
wGGKDXS0whywj+JHQa5njFEEw7VZqoJu3MC9BiWT0hcZWEge0AY5rUS/MD4GOOlXlGCtecGbpY14
Wf19VC30y9UgW/FARFJEoCmwHhQVMGfj8lVuGKrU3WOgFlXMp/fwo1K4HnV3ATOsj5qAIw4WrPgr
gwcinyM/MG7uYfcslQLXVOQ/sReO9bmpEcmlieTWvfXRJ4mM70PwY/xl5y8TsxpDaAg2cdKMrpgP
2O/n172TC7zbrl03dpk7emxKS8P4FMaRxaFdpGLKKtNcW7EeScGNoqYCvffMjL/ul1mBA2fCXqUw
DLCmeVOjxICG8R/u9wItSmHiAujvviOKI1iwPlTVTJoQZO2elWMU6RTU7omO9cnftNo3I4mHuRxu
Wb5fty8zwjfPcD0dstbHMVb8+r8OM7gh/bAhBksQ1QVPfc1D/G+wK063fPoJCsIcl5C/Eyick4Yw
NNilxRfrxjwdGYJ+T/FiyXZlySYJb5Vu446wi6+6jv7eRHmoouIBorlTO6EFZvam3FsqwlA5jLNM
OCDviT4Ag3D5QHOobEkViZr/A3tquQZM5dHVyHTXcM3SI7PZ9GwYHVrQZxXDqSWuZtnHUOnGtuPE
EuUgeJ7InxKAg2+5gbG9sslFU7UAFMwV17eL0rjd/TGf3o+jhomU9P5ju1pbcZKGkg13J9sjeUi2
KOWz/ZwLcD/PrgGy8gRXCttokOaVOSlKQwSzGovaKv1IqcpWKnkkMjwaJvn3ifzSbOcsabogzbJn
AVLDSiYw5Z7Y0qsc8bCAYEmEy/iTYLww5cg7epoc0BivvcfYxWJV3u2Qjp/WqKvkh+sSxioPq5qW
F0f6AxVzKp9sDOSo5dvABWQSEDdFINtfJjf1hBVpIKLmMDWyKfQVsBKJuo/umHqbShG72e7/yLnL
b7wu2MuCURtCUrkDHloOAKLgM1Gwm1AGGonNePw00IB6WatPCBj0JNSDEID5odJe/+ST3cApQHY2
Dh+JLOO79a1IKlqR3jSUpnjLpqlxL2kvEvL0xV7gvCbLrRPmTLY42CrRTR6C2QJpp86Senzmn4Dh
8hdufy+4oZTycikDVBcSnoDFy7rzHOREJ0d2v4a3MXprHKJEEyekwbb50Z/2OG0vzxaAydV1ZpAR
kiC9NgmThfYxEpqxk4UaGkaUURjri6/Re85i6Big1dhXW5c9Fj361Ig+DjU7jEuDw7v59ZYoa9fD
WolyK0dZPF0eZCHgjbCLuqPWZDrg/Kwb0LlXK6kvd1kC6OqqDIul6NCK6FWvpzzdoluZOpZ9g+kM
mYLtqJmtE6ZEhzo/OzVSYcAX0WG7V2WqwFaMs/suOt0y3JKw780ppkvHTViwkQtrCUiqERZkKPdM
NcnMSKRYueQYvMTcoVLMkk9iDWRrVhkpCIukY2n9iiOwYioo3RRECNlUz4+MzcUuPpJVRv/+B9VG
G6fllXuHvCGZkPipXTWvQODkft1vPCaeNjXJ0EP0MtfLRExV2W5c5+WHqL/q0CkOQmym0O/NYxg1
t1InjooIeG0a8LQCGZEfIRSfUxSmxovv2w4C7Hi4k7z5Bu9YQYXrOAmgV21xj6GZNULxiXr/beTH
o3CPZdv8XAlYhp0WlG7Dsqo5wuqKjTz7NKBziqWfff7N92GpMQuYDtSurptW/fzmZWWhqNTb/MTl
4CQs01mOq+Cyf4dbOq7IWykwg51xymaqcG+8bphD4JGzxo3sanIW1wcjzHXfMn5ByxJryqtCBxMp
/V0yJCo4brtYfbOAi5ltouHwhk0r94kOyHi8E4NPE8BlYWTAeTqsUYz/G6UbigtlnghGWANZbnwo
TRztAYcwIseGoO/TpUPFcvPhZTGUSeypZulP16ayvValzHdXaoZVBnzbq8UJ8KycaUm9bpHWyc9P
KCczZFX2Gi7NWQyhze7JWzuEpPML/pfa0tTQzzeIgFNwszeSgFzaUUkBs6GKaRNlSIqZhwJTBJXY
dR4DIdeyuG5/vkSqvap67bgQbKmQjqm9hNOp7ad7u/95rEoN8vdQHDfx74qlg/zhe5Es/8pk2kck
ayk5vr3xUnZJ6+IkvupPpKNQDjvREIpZwTX03xj6UnXmTDy+RZjEvlDbDcCssDwNfAl8hx9TbBsg
1dOVuC/43xxeH0Ct2GHNeLKh0XDzoKNra5hZ4smxN5Hdar42IeFN8FNTuHa700JFJXYAcqacX6+f
H9InkuQvwFMhcaYG2ampfOe+EjE2yOFXzdInSaHA9u6/WSo2KnInksHTuHrdHMaJTB9EsH37l6Nu
P/cN9wFiQn6huGoZ1rjfwtjGD2oV0/jGQ8oezDxX807Xmj4Grhl9k8u2iRDIsAOO+SwqBw2R38oC
8yl7FiZ6fhCyuFqQx59cjykJJKwkHMjjr0XWBKjNaDsPi2y1Qaa95eqabRNm5dWLV5NTWwDBVbqD
fupIGyrD1GGB7XhOpQMxAFLZA/bbRezMrM9mX2ZnbEYfLuR4CQi+NnLcesTIKpe77prToEkKwLiz
TlJxDrHs2+JHZoZjlVTNzrBFJjP6JyF0igwMzGfvK21cTomzs+Cj7fgqigM1s/jtKOeU+tH/u4xJ
guG1RbZKHplbXy4KtLL2G4RRvKgvgnVrtmEd3tWdM0FKr2elvntuGgAj1q5rbqLM5AKkLh/Gxo/l
S9sMWSKnedRtuNM314UFjSzAr4jHpgqkZGa6jpdZGOcwFw4p2KyAGauGCzwmPnOOHcYfhQNCP/Su
gIj154fsB66FMBPHWaxXLT0/AnJqfWtPK/wjSM+liO9H+s3ZePtPrCL4vl3CEoLvSyUuWkAtd0Iu
9clsOdwFHYm0iF2wHDWGvLQQFxdZuNcA7JcO9CX6GAW0QH1ezK5eoMZJYINQRBFRz1xezS21ql4h
wod689eYDsVTc8LzUk1WGX78EA1avUuXcFt911fVZ6pw/1S0HElgl8Bq8GziDtVhFXvPebdP64F2
aOM4FWmI+InMHMTpoK1AY+XnPRn1KlzBf2VBYmvslDPDL8T6zt/zkwDerJsylaKRfCglIWOUNvRY
GuCYT7NgwcrlwIY2nEUdnOiQzpq0Bjx079xNWzJskouOpXG4aIyPNGuhhv5JY+tF48IpqV+en7Y6
ACoJsP1wIsLDWW7+BcPsyOtC1DelvvT9DwX++aTpMskIs4jpA430SiIR3ggV5H59hsyT+0zEXzAZ
jl/e7FBDMlDKrd2zdZeYsyjXUDVeA/ts39DQ9Nj4XRmZ0tUFYh5nHhIjIFgksMt6TQvEyRvs8OoX
eigqj6v8nvsXTKd321FETGXfyWVCEQksB1I8Pmj6bNeEM539Q6Y1p6L9bFE4MEmIi+4SeXBI+QCy
kaHyM47m+HIq4cwZA+830xM8O4xGY3LGtGyYGVLjED+2QNaow4ZZ5+Xy809i94NQUb6fy4Lkk5ML
MvR3Y/68bjIt5fsKiZVXlowvaZGmlWoQokIXGLefzAcDGoVL7uvj9BcDv1NQ4b0NbsSfnDgTnHIt
GQlUi1a1znHrHA+iNVqHGqr0cAdr2+bpF4LS0cx5kd1pIYsLDhJ1F4yp02EsdHiAd7QLCzHty8Dw
qJcRLpjgeH2Hmv37P22BCpqHyqa+mmcHaXow6aC4Uk1K/GML79g3Mk4SOzCjU7wF7wrXyfX6ckJg
j9wq+Qmjmfvrd9hWvyZR9UqckNnX79eLNXsF2KhOGxd2uJEme30FMWrQ3Prq/YvPEBBzQuUqJqBP
1lTkTj/KKyaFs5oAfI5DivSpjdR02vCNvRZeW9HQ/5NlUcngC2017g6K7LNLN8DHNLscmyeRUsIo
yQJgek8g4YQoyjreGLHE5RISK9C/8F4aLmsy+RafayF03X6AwjqBV1ZQYJzWtqFR6Snhw/SlHz6Q
M8SF+pCLhR8CBnFN3RV+y8q8TaTG344IXanWd2EY0A7tknb28Od8IrCMOl0IGAEva9SMyycdWUDT
1SiOdAvfx/ZsOVcwxddHRIF559h077Y1Gsg4qBjn/SpT6b3bPxqnvGIGyu++iB1BXkHgopz6xXq8
lh42DBXQIlMwHBcHIKHhka/RaK3CCGeNwejdlpCxIKMmBp9ftNiVYoc/Vj0qYTLh8itrDh64XXR8
VQUIzsikONf3YCFPi2xCwqjnhtQFbMNPGmH8L/u7EMF54swwu2iLuAKK9RUrKxuZgKwjUdSsosKt
qpot/EdH5kvADRXWgRN2g+A84NCbPDEY4bzxe3ybKG8hibB5RETJIGjgDQd9Ke1CpAa4PBdmxJxU
y4EyO8qTo9VQUCCfcGHrI8pWN7VirM7ImmVciKTxuOkAsCZr39Klzek338fHY9zPxeUI3uAOgsop
G6BEjkBJfdhy9F08Gr3YP01NHNGroSTyW20FHwH7aQhlWu/mmF8QLAkoSU9jb6h8C3c73zi0qHUw
mdMB1D8ECsssoCqt+HPLyQUbwgrct6YYBixZYQdeHZZYq2UswZDFJSNIQQm8H+J+8u08klIP3Hty
Xme9I6w8FEgTkd0ITKfNGUHo7Ty2AvPXm/tqygG7+4/NWW84RQoxNkkvfBH1VVOn82B4y4qtTGjL
Ue7tLzbAbeKXvTmMjHVJlTCpmZccKAWqk2+i8Duwr59+Lu57QU/cGo+rGZVH6Zq687tFqg/2l/DP
WavTDoJwmdX67JCh7KWplXpbENWyVJBorJ+gB0oOPGisWNQ9Xv4eRZCr5XdnqMbkF9MwK5zCMjPn
CTrRz1wqZCBzsj2Tkrs3LmHv2w2SRpo8Czy7z5QUS2fCRJqlJ3hkGuN9NwKlLaL/hNk31cRA5s1S
8wSK3LvryaDd1wrNIWhD7/KihmhwuasBmu/CpvjHSDxt9L7GPekjQ/JigyfeheSEN5MOVOPyzmZ1
YxkhZdl0xZUa56/v8eUdRoV9L7ZORnKbe4qzAwaz+dBZsIYzt6mpDOki5ZYDePDolq1ZnIo/oWsB
Q1jTpufJScjdEZmL8aJsuwB3/my6atC5z9H057fRL062tpq+zXhldeMO2Amurib41pt4zzad5r0a
Tuo8G2tx9vhpfgiE76LU3BQ3AF058lLTVGMQNnN9H9l7qB5RyLQgiQnR7WiC/drFStDqYae0A+vF
wbNe2CAindHin25vxQP8nMkJXFJB7W5RG6XlV3VT+vGw3Rrj2hS1LkCxs0qodZKf0kTmtM1r6OIU
1zA69BZfqz3u+lF/Idy3Se3MWsh4CodktemO8UE2pctqpacxUX6GyMnismV3yqxibepgraQXmf72
i/A7aio2ePrMdAMbtf43MJc43MjjhEtNAzrpWVvbvWruYSL38TaTqFKpI+gOsnhWu/vGmXw+vD38
Uc3J8wBRq4O3JA8yOSvcVKsLgZxTOOrHj6FFkCdefXZygEjrewZgBNL2kSaz15Sk52d8aVvjHoLP
eeAuU0lStahfDeMdaeuC3djmdHv44qOij142jJwqnVzHmDxYW2jRaYFYFEskAshvRKiB3kh/+MOl
SOjBqKprI7fFQQpIyzoNSwvlRh0hnQUHz/Aux76xiMu+9l97BiXUZv7Vtxcuv9d6UhG0CZzSuuj0
Xqfn9xLIvymjrGGGODUazhDVX8RM5eWiEgtriSNPKWV0bXcBlmOQSL/0kVMJrK6tOFJTEopQR1co
8tmEygXgCDI3lvuxgrB6fxxmgsGbCq82KZXtgJA3IdSFR3JyATJehFUvxV6zGfQfGBRrVE+HOM/P
JuiwQ9Y8lcwxDitkd3DKYq1boEcruTTquCx/seh4zU8UKsq4cLzCor8zyhDZbeBWhWOgTMRlYY9r
86+oo2I/ejCcGc7xDTzHMvpQ1Z5tezn2dXTK24+DY/02HpULQH1ioPMZ2bak5l9gYz4UmUjusNrj
lsXkmWZdmoAzDg9Gbfpk5l8tYujPk5/Qz1loPtlbn2919x8i4c1AHfQbV2CNTaojzng8QVapIgys
Xr23MnRiSCnMTh/kGqFQKgRbjW9mXOv3QbziTSf3ScSlLqrJ2qGdmFBdVze9ZJeD5dNJ44aj4ESa
7HZ+bO/mSwzW0seK+TtdOxqqw8cX9uuRGwBGuE7CCF1Efj1MMsIOI7lyAqadjRAMvUquKtWL4xit
JpyYCs2fi7Q6Feg6xRr6hiSulaBncGZ+P0OgFz0LK9PCkWbVBcH/N1ZUI9OxcWmdf56fGbitN8eA
p3+HE+mHBH/KcRaee3yQwaCZeorOPbL6XVq+5w2YmO/HRRxBvSix51pTJcq/p/gAa1HvdW6Nstog
S4yIMLvt2ozoNvPRPmbPP+Dsvpp04ssnKCRNEoq6hm7L8C9xqh/KVRs52nyvdW21oVnzHabcF74r
i/Hw/+ssRreB1IpWitH3RUm//tLD7RSCkhKHWTIv3WKfzkP5Ax8KJKcYNslAyrWAyM0p1ysa2tnJ
7zXsYWHt1jIct70af408YEaES4AIIyHVmNdqfIOnJoFlbId3QDG2ha5whUboDtbtiDsZwBBMkHyL
8cObAvccVmDDcE/IxsvLjHvttgiF/lhThsSG8fMH/Nz819Tjr8hrTrwO6AugpE342qYr/sH6JGW+
WJmC/f9zeKnhZ6NgWlARzlPYZJvHqfW/6yXtElH198hRa7U6QvuEWeRSjcX5KQe6msp2TemFrAfL
SALvMg4kqsPUlZFiYvrxkjNyj3GlNUK41wV8ZEoKcTee0u/jvwjfinjXXyF9eLFqKW3T+I0da2nt
IZETtgYZXq4lc5cUhKAUygkAxoAvzfQ0VQXZKKo+n2b532+n74hBeMpFLYPJifkdiA6NWPSekL9S
UfKybT6gfnE6B0ib5rdGGOINJgzO15uxqWuNTVjvCaN4Oa/eDcmiHTBIpNcSbS2jjIQbIfnjGBFf
1TnMlQzsaYZ8jDwzVT1nnXedVczn8C1jhPBkmX+OKQHxOKJaOLhwo6xORrNPmjpt3NESsEZq/ZHY
CH/DO0d42tkP4MNAkpr2G/xKfQ0XHe4SjvQBY27chHVCHbzpI8FsE4UxMgTQCdHfjqK3K4qls4dF
KidfuoszfnoyneVer/MVLwisyPYxuogzU0So59EVxEB8VXJus+Ph1iWV4b4ew62lL1QyaiS8uG/F
wZ8fI8GRkb0m8J23GeFD/wOkczSEhHUN8t5PjvlEQ67mlADIOazJB5I1XW+bVQFCpSHSPmjW8MSz
f8pTjFadK0baqtm0RL4rkV+JYdWILOF2VSaUWp/8qRVqMCY8x/q4tIiCrFwpqvSrNVP+yxhRJDk3
8U9xe+QJuZcLwLw2LLvRdkoRAo2rj+iLTyNxTqJ1DTNDUdfArdzGewZrxYPN4WyRzqvb4ifu7mui
xph2q/3IeT/CkH1g+fazLUg7Tu5N4A0XMbbBAw7lercs66uPoMtk6isAbRo7r6ROUQ0UJPvB0n+x
aCRWJ82SxYyZE2h+CRoV03t1sVpVQdPuS98HHVLOa6yB+kJQ81HxCpBNYLwHl1qFjHjRiouKPFPQ
z05vgFAtMgkRn7Fhqxi2/KvmgNZGkBusRHdh0cDBcTOTyBAQIcwhihrXCCByUAX8LHrebaxdy50N
igVzPiwO8HKH4pEjfXKUZ+QCzKIP0G8odWe3amO96okuFwvMDazO0BVP3JHhI8R0OTXeCD/INRNz
DWirKaOY/09Ad+MVXa6vQIXWWktjp/Wb9ddXUGKzR3YBlQTV5peLbEC8HCzq2j2+BjRMJpd3AnRv
/1hxemwUp3nyfmEvf7lMpS7p1UGP+k+TsqM9dBDA9zhQGtznLGQrRFwTvXrXU/DGMru77pEFWh7i
jeRxQN1ACbSNJ05qo7gPCLuz7ETO1ddqpv2ndqTucnMWwqMqujXcBpjJv0sxhXRbs9vNMtVXLdEC
pfrjckT3zBhVhOjK2PD/gCWSB1RLeqmWKZZfEe59PyqP5T+tGQSInBF5EyjEpHUG7OZOu8Wk4cEs
TTulIE0NePeZQln2MNsvwY3THBHz/eSIdQlnx1otxqEPlRKvGaK2t7WZc4MKHQxzScsFBThgBkWO
5d5yO3p4MohddAZA+xvUBMDJpBd++A3Cm4OrWztOtA9gXrBparkBQqKWk0Dj4b1wZe6AqTyOaNey
FpvfFOWCJcrciVzbGxMAXgTPLy8h4TixZiuQfac69aJJeQfPdScfvlpVWFw5h9gXsz3hsulKWUr3
/NJy0Z2h5fgxeevOCoGwKojxI5c86VmuxdAHLVrW+6Non9n/8D0dvqlkM9cyf3oD0K/wno77d+VV
pwxdaXBfyD7qkBoTWTN5mcUvXHL44p6J+58ICrrbXwEewljaajEUOvO88s5df+vuvEK1lV2k2q60
pTDaYZu8FjEQs1oJ0fxYKupEWz3iEx0QDEdTSarjeWs/nLczTQB6wnh8zKLQIWBv5NCXU2XSAPYG
zzbByd5Gf1g0C7vVOgCl2DWqM8ZZLT0DJjETpysmfrBz33jFPET4geSBciGnVPL0HTWfu+OQaCdC
X7KjTMWms8hvkuqZdXnfc0hrkHIdtX/tHGBNygi0FKheU6OhTlsbkKNrRh7A5aslp7PJuLUEA6cV
xpe7dZa2AJ9C0GxzIWfKghYY2C25Il8RnbiezC/QAmt4XruD2O//2prhWUh9RfZQ/CKmXMn3bCZd
9T0Vc6gUJoweWu6gwoJjHtyTGMh9dK0gr0Zh1nn4WY+5OwxB3ZKcFAA8O2lEXTVSpsrfhYg+OXzr
svPQr5YM7AHetDSr1eNnOjmo5DmknJdbjDv185dNGqK68Yp1xkNNxBJCwErHLNuGEr/+8mxpdyFt
2TTyu8iMOPYCmKV1SGcn3mcnwAPXuLcx2wKdts67Qm20FFKpoBV9mwv878VBYuTBeD2lfpO7/UZX
ixKxevIFnMF2ZvMDKKnYN9JNZ3ZO/CjCcuVbOQ7OhUkMdL9ZsXZqPdLZI2l9jPjlbyOZmMzstqTN
l+F4+TJ7SNGOdc7MDtFEg9Yxyx2XbAYoUnhlLeKFY3VwDzlOQFOjkeFKLdedMI/cp21lznmlSLle
FDsUWcWQ2EXz/LvO1AgoIYXdrIFkCCRWloIeFUi9Ojok3boQtQX+9pwMu41Ci75yqC0WKfYY20Cb
F4fqKTa1Dl/Iq8DOrJyNnbp4O90x5OtaFqtbtRgqvAbOMFbxQQ0vd4b4iqOb1L/lP1TM5zgb6aWX
cwpiibvxz6nsQxi3SlKP2v0MIbpqx050zK45lB7QDmNspjuRBH9TRW6KPMlbCxyIv2acIdu4yqKD
7TzXRdQFWYQ6zUr7DAQbwE1eXK/9uEiHO19kUpXpDpNnSorjbN2gKPaqnTal5MsHv2s8iAqXV0iE
fyXJcdOTJLrDuhUdsmKOmvmU+0g8tynM0KOSlzJQL+WoLN3oXQpFGKgBILZaw8onJjSYcnoUnenZ
kLNpEnkf0t7n3E+lf0bNQkLQaRbgkwl2uACUo2FfskwQfd84PyJxjGB1ZJdeQ89WWy9UFNSMzVJg
qpT8c/ULXMsDiOG5LfexDIjlbP4vBWe3Td8OtIfSKrfmd89IJ12fM3iHrJHAUwZvfVCLx0XwYQtQ
wdg+pu5oxQSjFKwQWvz0dnJg8RGBMesQv27sRXbFm8JNJ2F5gEwo7IZM4xSTDZi4NNhu5tjMBmQL
Jo3klNA0W+ZGBpvqd3u3g5mBypFaVWXpcSLygueamMLpzScTsgyNs3gG1pp+eN2F4DnCoi71vao1
ECiX4larpkkhxsnOVHcrHCKSg/MqDd7vdd4/tq6zWc9nw6iXEXpExBsZJw57mgaUMU3K7rpQ5hd2
J6/PK873IIOVsW+4ctpl6CEHjJGXCLwp/1J4ggsYPV/zoMgaJQRfjNVKfVkHEC6shA6YZBxZJgON
goCzagtD8T8l9niXv9BkJmmYjYcEz/nJV1DZqPlsqQXphx3FGB2nDsqFlmgeLzk+OCuFyQTa585z
HhDohLqEwEzFbVZNQClsp824RVKi7WqQ+uz4i2wXTzm4csKspT7T/LaCNb6utyXvaeacqIyfd69R
VkfWZRCKiM/x2bJFodae5aK9QMxYoDH2jejL7bqAxQQ92HxyRXzPNHOTbmN0VBxLoK6V3Qdv4RXn
F2Ev3LoM75vXtz2cCIpEOiELNGMwajX8aqQr0oARiKvbrm/WehC0uSiiq2gAit8q3CRXDKuh3uJX
mR+HJOyu/SD1ZHbTcexWTr3T256oBnhjJz5ryftW35CZR3JfhQXWtUC6tnPZF5Jw2jlcBw5JdNzR
rA4zatmASM6/F9mn+PYt73V5aoFhx6Aw6IXImMBDKLuriib7QUrH+dJ/KyBLl1am6GzKhLYyTuj3
QdIwk1XXuqQT/jVcLCzRz0Tjvr82rstFofIpeC968etJcDvjlzdj3r/ObhXVNAclBIUTgHUc4V88
zk2WU4HPoLWWl1SZphG7KyZgr7h9iyFEH8T0ZHDx3V8CQzlLgMmINpg47KdP/R2p3ftpLfbRwUrn
DI8JluUJdM/gmc7vVe0qCcj7LERzNU68dxlSnqIdvqJfU9AwzeiIg24lRnXfBSukc9+BqL/v6CKO
y/xXs4mMH9nNASAlMQwZQ2xLgqqnb/zZAEvT3w+jfrK2e2aNQfal/CNK0PB+mNZF3yxaRZvARi6t
0mDU0C2gWyBDRQB2zSRDyPeurDpFUUQJVh1bSLcyU+Z8Fj2YVzWOgeWd8auOgTO1tPkMsZDv1iWD
26W6BSpnkQ6fRqnl0BCTIxULEQo5zgTpsKiQbRU8lZEX5JNLFgtLJZEoXD6o+npSs8h5cA9o5I8l
NCKX+h5AbimpChNiJ/kJYETg4XORvwa1N7iL1SeVT2tyVAk+OmlkKcz/YEOwtSodh2vSkX52Uquz
sc4LZziRb+fkb9TAuGcE2VsLEwy0z7qz1L3n7zt8D3n01EBw7V6R1kB/PjLShT4YXRNKVa0QMTho
fEnLNIiqngydVsYF8hm0l4gwC1gabzmZlz4pW8GZ9JpNFz42eVYj+JlCaqywE49ulYbWABdLv36o
lyIc1cx5sR0uvZwVxIG2EBhOYbZln2bkJZkRVOPGWnUuwkVNjeQAaguvC5ONWga/1mnAWVqnWUBy
L0FhYjgDj5I10MkcDeF0BZah1QYeCE21N1PUXRZk5Am8eiPSKXhNfWTMuSuC1h5c1t+JS0ICsW3A
DffmiUmFg/fhQNavTrTcW5Njww4matZSiTGK6tHNfTjKnnE+pIan7LU5wI5W2eKC8PliGQu/APeN
yliTIINwFYR38VkDMloJVtwufSs/WjBFRaQ4v0kHPEUOpcKI7K+FA8wlm0X/OqYzUx5ohGeOtQbN
Oyjro2IjSfClQR9NEoszxBC9zlqlzK1N+cdDAFq6Mar6vfJFlyPsx10VxUYiuxBIzDT77WrW//Lx
gP0M71W3PYDmSY67KB666pG5yblnqk94gVSmWAI7+AytAqlr9Sw9ZKa1G6COkrIXELhTJ4o2RmHX
KM42i08FSs2kQo9Y3in6RzgVNhcKHAmd/s0SZlh44nbvpIC3ew9eoALIYHGu28RU90nE2p+ND8Ya
sV0Gd+TrzteWPd52u6YpNU5s5cJ1HAwm8KxRwO3v7cz7OzYlU9SGna8fNtGSxqwCl5af5JmmzIow
gqkLyZL7HR9iWAER2KN86zDeO1cgC8VHVJn8Hdn5l8wtbcPgc//7hXW/4ri3cuBUqDsWgpX8oXdB
4J/pjlM8cIAScvx/dfwAP9pJBaLIMmwII/JdhRHUnc2/Th/JgnxDF6SbIvbWCFfpF+xPy+AyjB7j
csk6z+7LItc8lvZdRwhHd6dukocx14BWd443ySNx08+GhIbVjYy/89EKLSC9mvEpB+TL3Uonbful
Yqswz5clpmodaaEqhLvCfsL12iCbyQ9UUos0yCEVjExRMQhiNncQ7Cf69ZisrHqUmwIwMMHKrOow
Khoc2f425MhGxcKktpd4Tgd9jlUDp4ugxeZrBRcaowL2A3BdNXHJn5lLkoaEJKlGGr/PmMF891Lq
BV2E+9dQ6uqKSKIbjYYvfoNsQ1KYgbARZ4OTaizamixkP2uW7KX2wrBNfF7fxfNtpEGgbAIqCoVV
gn9ohF+JpZbxtJFFldtuUjboeOJjFvPE1qCwr5q+wJBymbxBboKFOvaffWrBWX3B0Y+MhAq5cciP
IA+csDRgj/DZP7Wp++/DtPJ89xysJpn3Gu+nEGld2pEiUyT65cLVIWTyDfIBsOW7Ez3T9yayHLVQ
KxhUGBtSiGtmWOYBjnl7xFl1oPzakMhdiaIc23gTGiYHupvAn6WmX6VGjlLgnamBExRZxagBBU8O
5HgRR8J2fG8XrPotWmZWsMS0HY/3jml5CPuVE6T9Co68jflSJHdd25Wo/kwzeWm1ch/B2Ug8sjNI
fcYPiZpnIvdB1eYVcDrsdruU0uE/5MhZ9s2SbaL9kVAiw9erGMRBfdB0X3SAKAzdMBE8+ZVR+I+1
50Aj4rOHrPKtry12YKOhAzUDhw4rb3e2x/80Vh/dlR5fAK6OGEHWZMMUdOq+76J0zWtxBN5RUBOa
G72YlmlX5aHaKgOj82BtrKJcFzpCajY7QuuqjGuuNm1I/FRrh3o/l0H058maYPTk82ySf8I/oMmL
VXpUpq7NPkhf7NWWbiRMyfUaeaEOni/P5R6wgYvFxdF6yK6AzBDurYPD4yWJWk4xkce34U5IPEml
9S4cLYe7fgtDv/izPrB9YEyL/YLk2Dt83UsRqAjyLpp1RlQBJRnk/XffbQV3owOnLlKFIQUPFNsC
BMLDtzMeN7mAJtyMhzU5m+McRWKa1lp36/SGeF79mYM3+nVS3nFJZm8By6DNV6GZI7P8htXu6Vty
oHuZxvOdTrCorzT2/xWTAd6oLDYOiAQo6LoPJwTIjJSBA+H8pCQD+XSBjQkcDywIsSGhRNOCycBJ
wkoavft5VHIRu1t7ITW8WyxrfWNEtkuy0jno5B4AkAtLp+X/Rh4U+CXq3dvGpZwxaRYdQdvxoMKL
LOrU+FOjhpuh3igjx2QkG7ap6bBMGcHplN1fEsI7wo8gFhuFh0CcExDR0I9msPjPxIriSpZLjpJe
Jq2BMJCNanBznh7QeV2f7hiMAG+6JKBbaqpjqyEqHb9h9+fa5MgWb0QVQrcfxu9pP+9phlxQSwpk
p2pvgbRtPfMC88a3fJn5PYhQSmzsGTwHmJOxFmOYSeJj0hZDobanh25XRv23GSuNjWMBCR2yJfQN
y9mAbTJJKAihNIXk89+kNeBG10NZr8gIBGcafvvYz5APVXZ9exbfSErdPYzFP2o1LOqQJpnLjlep
7c0kUDwFs2SuptIqO+97odtES4syA8Fsr9iuoLVKZoHIMfJSL09JmXpLJzydfDR8neHjpgxS8c/7
M0OXB1eXbqArsW4OVIKV9aC5tLjrXjeMKAGFUZvMFqTWGKsIUK1CyawIkeRWiUjMTgH633k8kuQo
/2x8NyyBeyzdApBclqRAEq4IMimp//U9JXDmC4hqsf4zLd+U+Vdl8w1M4WID/D7rzxHP/y8A1H8g
PPxYjRONj7eCLeu/QVLXy+R8vMzv4Xfo5Z7aRnI5dLBititgnGrCtaEAK4OHukun7Z8q7+ax2GBt
9apoi0flyx0+SwUUILj05wwG4/j2oQRbVaz95OwTryE4uoigDeKWWEu0UpgY863sM973d2gDEX1K
pkOPbgqIYtWu2t9ir6a5QHcQGUHoC24fKCMYJYeYf57Juy8g8QmihtnbN+u14BEubrh34v/LE4vY
TMwQOzb5nrVlSCkZcMyaBHqRvVBN10zlMAS8HKioy9T4M+O7QiBiwLp+KBETngG4UOwMwqafRSLH
Kbn/lAk3mcybvuxSa1tv5XUC7DtqyxDJxajuEMLq8aUiJ16z53vym3/fX/65T0dYo519xWK63x/u
lE5a0ZbCbMsa2XH6PbMQsOT8jXaFGxy82VppURYZWwAe3SAjvHP2sumgdYM0iQECyljaQZPWRqQL
v1kB6ln5j8PcwxemlCL94GSDOW2hqKPicODymdHJ6MllBQ2w7a/nRxqNFp6zNL0RLSalRRltwz9t
fJ2YMEdllE4uvMXRFDFH70s2bd3iKjsxV0nNX1je5b7ejQ4MqDoz39DqinRAjNaYBuklA4WN4j6z
Tlz73k9r9B/8wdTVgMa+ju+bJkzkL7Y30B+UVBmMNyhAJAcVIdBLgKWTv2b5o9HYC0dTkjrZTXAM
5goV2v/pqBVLw14s9huX0n4vodS1KjwlC+Sv6uQTWHEkB+XUiL6Vm6wR+iv0bSGYe+K6Q/ei5WPW
59s8cqi6stXzAcULgc7OVLrewZSuYFdW7E5UnV2a9NAWNk9HFpooc4WjQUTVgl08zqeHnR8GFUNH
fVnM3QNlMsPOcs8/AJs6ZO0bBm86f/lJHhEwZhRBI4GN6sbNunHoLfpOxAVJTwMfBYOwfkrVb58x
5LaSTHemgEU3OqQhopoY5DaRtY28xs6tgmlbAsYcoyFm043dBcvPWVLQdNUukMoqv5FpclS3ujaw
gWykooThujuMca6gdW2QbLdFnJGeWckwBpjwqUXQFH9aZ6DiAHuSP7aTPExbv+ouizKbH799xBk7
yDoH327vBDjCX8VqZejeJOfEAGCL2m+MiHgE+946xl/SGxDp7/h8lDJ14c6hWBczZbIaolZF2/Md
joSmd83T2eSBsD02YcneInp5Pylq+hp+Knj15YZVdf4k3ztQEEAguI5uI3fV16fHQJUG46hC49yw
n9FQHWv3Vd8G/dyAVxuyxoxIRy25FmYwA7WoYtWCvRME4hWa5v6zwFSEWoMbhhhwnkO8pR7aR6Mm
l6eci5Noro9N/+NbDt1WmYWK92rEwtX2F75g+WUgJW7fmmCWwEG5eGBC/QKR5lkci2Y/eDwGfc6L
5bc5QeWXD7q96A30nvYUjhqn1Fog6aflAxNouAxIFd9q1HtoCyumG/g6o36i/sp4s2uH2rUQR7Lc
0Vp9Ms2Y7g6VNeT2Vo4oX9awPn7ehE/p1ZhNVZwTVPRaoTBJtyzy+0J4HZeu1DKR8Lx2b1T+xjOd
BQyEF2aTIQ5UE7Tt1ptpF8aTZEor6VuHI4P2ZWReNdnqaiDoQbpW0UgCYpEpkdz3w9XX32z/ReRu
fSIRz/GRTPUTKt7wrHyeXclCZMtVlM8EjPCN1JF/wRXKujcSLMsp1ns2oiuUENhlZlMTPbjs1pOL
5IG+G0lhRqKYtvUhHctyycTsPXsj8aS1+uvPac9/MayD6IzIEJ4ITSEEO1wXMT+aytp6AXbzmmYW
HIgCTvXAaOcqP84R18MywfGbZjLu+w6sExZLuQhaAJ4rOP668np09XkZjwlafHsQs7+Z8mfHiuU2
ssju6vnaf8s7xpWc4cYbBwDNOIzV3RR8inDD3XJU/oSW6PJOTdAYh3Hj/lz14AU1I+D7hdmDFyeU
G+653TUJzkiRN/Ag/nWTYhpmyekK9joIAXYPtcR4A81vEidBbJ40zS0n7WKohIyGyfwfm6kpEtFf
YJHTaYIhcyOBSckAP/aGIm+EE5yKUxD7VTqGcmncZwnHu0MHX0paAo8CWS0J6MZMmRiPX5ghk9Ym
1N3nTb7hMSPVIIMWt4bbRSFy+IN590oSNnlU6g3JdmGE4Q1qvSPa6v/V4P+rN0ur8c+xnkBROSLy
TQ412H0RZbwhvuzwYwhWqA2zYMP/ndiqKq+n1OLihD4KDzs5nsniKYKUAkhkwUBZeBc5vmg5e9Yb
DBOgRzekRIiKGWDim45o8KhrS4PM3miucOX0RGSx9KKF0aGGFG6t0kBHjwybq2PYrMepRsC4cIvG
NqOQU7MaOe1Mn7K4A3qn5nkaXlLUjEczlz+Sx/q3oX3iu+q6b7HxY63O3czafnegDGhE7DIM6YrT
/jYQFH9CqF2B6aJCjf5xUG9mafQGeC6C7n8dbp0akJ004Zm7k3r2rIgdAC1FddwmZsOgBYyakmj7
IGJDuzYFKFmA9Cyfbmg1y4tGbe9Zo2TIS4N70qd4lYFWV4HlSglsWyPU4pT3VNdED7qvin2Cz5H9
vp6Bzn9oUoneTgI4nQvL1jrP2ZE1Zij49auJvj0Uky4MRCTMzjnzwuR1MBweJLQUEmLG23Co6Flt
Oq0ZEmmihttYnySh1exmoyCglwaw2HPTCBjzFfapk5DYJ/FQB9hyzOdTpTh00OzhCCukHupemaKb
MVuiEZQ/zDuBvh1BJc7O7KVXwaHIROZ5GKrAyaWLwR9/lpa2xfugCWSfmtFjXOKYbd57tZ6PbCXg
5mFTR+rWX0uGtRsfGIEuwcuSW1Xas0ktuIlj3oFvmfwBw6coCg98VC7p4/HfXTbhc5t04kkXGXjB
0uMajqh3YfTit8SecUL7cK07pBYxXIxsKaxMEgDxmUPnnaZKZZs64PGDxB6PoV93owbu7cweXBIx
K9OM86tN/Ca1+awjkE8qXAxLvmdfVXbbqTlJZNLCPt5zjmOFnsfR8GMjutVBh84gthNJLRXzZmwS
E9SseVjzLy/tt4QD0ZYbc7Ne9DjkQ7gM/ANohHDi5NJE8lmIKiX1C6wCGZcalnJeR/2ukAAieYCo
Z0z7LKAH3STzQ7wMmjS2Gj8NC/2GofI3unlW0FcZdr1OQY4Fg1lxMnFhxL9QQn85jm88cyEMxec6
5t2aDTECKyckeHnffxxJEqOOA6Za28yWe4yRkv8SWrbW4+WL+MnfpQfikxkopb1F+0syJiuiJbW8
/Lbd0i2hMZD9fTyhIfS89eJsqbBzU/ZmzJxMeGtQP7TlKZhDxkk31rbBtkhaB9YfXahfFM3Yp5JZ
/NE2ux1iBlwgFg3IZZ/68y0ri2t7L9lWBhuV+yInQe/7G3txMbTcx43/3hCnI30UAcLu5bS+2a34
+0IA0L74SPKSNnqZRgeejoNCe/XphHjdaNqH616Q9cRfBHwRT+H9W6VIM7Y00pTuOQUkIYTspXIs
HNhuNH5+5zoIdHvUII6X0WwL9donjvrYv7Dp7dN8I3jdv+fUROwTjM5bWluuK7nwLzhdyJ3SBBT+
zFmwhmmeEwBgaJvnGVaL+hlPvN5FOJR/nkEwPBmdKNnAnNWYCj3ZypEG/nUpvnVLpykbliTqw4k3
qWNvwzyJZDdv0DXzXQ1lJVO4OdbIMqTIwKsMEaYuVGG8c+H7W/wR8xucb/B//kgrc2WIfU246fJT
coqpdi9sLPQZVaOBbZqYE7ulytAJpqB0h1wL43YBPG2U2uxxVDO1B9lW7RjG2u944BJocDCaIXo/
SX4I/UKMIIsEvX04OcTM0yDkCuKio50sPUCz7obngBV7jxOGecVSFtc3xN62GO1phGessYqfR9tW
OazhBDQWiZEVfZf67TI8Y+bH1PypyXVoFHZEIsQq7wX/VcM1UVCwiwTDGWcYz+CiQ1LtwElXbmwi
WnBAs4fnOmS16pD5xgINGqJp0d0nTrDUQ5g8pjWwm9cU3c0S9y8R6TSEqbBAQGYvLzuISSP3VhKJ
NdScyJLPzF2QWG++877/t9MKy+H08sJ0xhBt9K0CP3sm4qk3+co8rJZYKVoKrzz15Js4Qyt6gOij
fHFtiee6h/mQTS1UQInEQPx5T41FVAuGW/KF8CIg95oPZ/FaAyupgnVIw6DcSGSp1fL+x1Nuqbbk
u+m8C6Vd7HLlD36DNu7mvM0HO1CfPbDWHqFfK0B6pK4nLlpjh4UVggmlOuHWgbZjT0FIDJMJwvsM
vbzV+34Sl1/fxgi9CZGHDpDn3y75lw6y6vdIKiENDzBugS74q7JPD2SBpTGBjmdWytI7praUBHgl
/ebLUwWjWdMnVgI1V5fRjbGabbSkQUcQS11lvHDH8Totu8De/2dWZWcX4ZVxEcZriVqy1OOkygCJ
quWrZ6fJqXhnxJiLP9JRYIqJHzf4vb59ikbVjlqUMZ6z9Pv8CGwRnhbPeT6YkUFaB+RtV5BfXI7q
NB829devcRFQPD7J6QVg4rNuaEc0mRLlrLcxQLcFTiDT2KYVjkOapSa1mYGw01S13DDgBUQtpeYN
O5zr/VB/UUzOHOpcIBHCqk4YAAADYZeuEMpswd7HeRLzfI12JqRRsybcOCV6IQsyek35WAKwn8Iu
8ajMYkqx2NJIV6/2hu7RoYC6/jUMokHyCpnhZ8veDhoofqZcvm72Y9/WxYKJv7okqdv/zwkl3/ld
KQtVahqh241ZQ082l6pbc3xvwIPIG7IwH5kvxqZSIsy2+6/ERKBEpOCJRm+mFcppS9nFWQPJBZss
aorYGSkYpIDf/+tXkii9Y+BT6XJKzyBiel0RY84xWP52awe2AYiGQbKfhp/iLwf/xARvkECYdveO
+RcDw3OYQ5cwBKnWFcr43Uf5GaqwQRdcjmqZpQFk+MgtLEbRhSdgEEu0Yfn5kDp22va2Uf7FqmhB
UWUJuBd4zrirRMAbDT8nB25GWO+c9LVxFGthnmasigzkrkm7UqLnUEQQ3mtrXJVg8bYjLI79j4IL
pxkHBFXzSvSh7H/boRyAm1QS1jtfF7lgMB80oQFH8O1H7rYiAyX0UovQke7GTg19tLX6G7RegiQ4
tTrnH6Tmeo/GDMlBQ8xSHcwPGToO8NUKGUm5XZ2cVHatdMRo7W6GQHjPx7xlemLKiQIWSHdNe2Rd
9BfkjDiCmww35scdYwqrLSTLF3TQwQh6R3GGvE4cuuq/xvu1izdEMG9pKmBXAWIKdA+oqBFAojm8
2CFmYUiqXrzhcttfg0ls6JS7ltcGoqAmXne66Piijo3SpBYU2CrPoPvs/cJBYZ1Syyk5hGy7eiSO
VxwRK2key0BpvANRcMIWoxOaa+pUgIC9zstb6Osr4oqL2NIUxj3XY2oj8bduU4HLobdGogZw1Wuy
azKT+qmqeXcvyQn0EXRFoK6h8G7cQFegLRSWI89WUJzs0JLv/iYJGGpBRBxdS+K2x4nBoHR/0Jbj
LB8T/WTRDbxwirwWl2mz/7HWuqwFa+oM7sS0JsaaYWz9YhIgVPr3lvG/24c3XGRCrCStmVwZnpVZ
Fc1u3HiXqSswoWH+eqgda1gpLG/r00yx6k+ghUOL8lgNEhF7U/yoGg/5+OopYtE6EvPgatMPWdAE
O37yNFTaSw7W8NlDlZ4OWwAkSixPZ3iSIO6v7xa+mU3s0BQndrNLAOR63DjyBvrJ9SohIpAG5XBy
MSZ88BZkif25+2KUdKBAcTaEqKKhVYd5fwRENfQONAl7kBksnGeCpT8eBbDBDp6sSuwWQ3jMimCZ
WI8MQFVdXN4H35YBWB1yUmLMiNHBAH68o4d9jJksl6o2NiilDmqbVHuJk6KKoYC+7diX3+XaGdTC
mcxgwBwKgzQAi0pbT3H2P9m0m6Yt+t4oDCaMZeyM47LGk0QRZdxKDZ9sXja97liL9SFTYouVZ62K
2SAF+DzTpZgLRsgMiis0HXnJmZ3zurNrJdaaZu8B0gmjeBJq3IBAko/yQndegZKW/XR9eKoXzG3t
KtW4zVGT0SeLoT98iWpx1MDkPhd+oAUqC+d7QcKECUi4Ih59MuEtqKmD1MytSX5Dp8n3Txp73Vpu
PpmLgDChKps+Fql9AK31Okn6+3PBk2PbTSaI2ZYhaMrIJRHbmqW/cleAQ+Yp8O1Bwd9xUpdu0uvK
wemMJNnpIKbHbytXBasK/c9k6gGusGFEqlg5f2eX7xCebGpHU5og3Qjm70dHykwsDiOtz/EJkKgy
icsgMYnhd8cWsU6Ez8g4Hqg7+XDivOxdkm3a5Ed6g2WHUp0onPqGxemgP1qwFHqNPGzn6PDLcxxZ
e94aGkBJIZUiAmI2ubosCu/McKHP/Uzdviy0xvWxXGs0Z4EGJLy5l1vA6UWIJ6C6auRTGprUoVAh
ilv11cI5vLh+FK77nHI18zlPCaH7sVY4Enmx/t0Dw12KgNotBb0PjKu2KAUwATMQadbdZuZSDBXX
OvaD5Q/T3LlPvaI/RZfg6WTEOKv9zxJJzuMQdcDzxVGIfncmfINAGa3PZ5+v7c81CVhqzyVMS+yZ
nLKHiUcE+l9d7GS7bJhtVjQhEcsB6/qdG4MT/yw/LaB4eNO3Ih5BiSNDXIkYznzfbhoTgHTaoJS7
GrrhRKzq4/fx1SshYF+mYYyOEztx31c45vHKZ8/o2JwpED5y6s3PsLJhRhVOBPZJNH47MZG2DMkx
5zrGYvVCU9ZKlfFqbfAUzyuYq45b3ZGvrkjS4UJeW0idEfNHWA4i2O04iP+Fz1x3xiJneniiGuoX
dYowIXnAYeeJOMNhFISzyFYOVwWq5FT0vGfiRw0QlnGpOrBH7de6IW0jQv+y4o8j99f8YcGH0tII
xSZU1yFieDAVRJvZQNWEztSIJjUEAsg9U1b79sFuprgN9BGf0C2XH8UL3aj3sgnjulClwrSsm3o7
AfonouYBKF89FVfXIdtCM/XJIX88so1xhUrQEezBvuikpXC9685tXSxAp9kl7pvCrp5zu7dt1DCA
leLkWYSG6yRfwpdSCLX5+M81NI4Ym9e4+M/II+0KLl5gkmntvoBqG4tL9Y9oPnPQv4oIIjMVix9Z
q1jEDLMkZs61wPALkv68IiYvTTHM7FQUr2ajbEgJTvo8uyVnRDu/pu8yka2aJ1OljbGxRNTo0fWU
67Me1K1J9sU/d0VgAndZL0qyPlzIDyYh5Tc65szqDEofSqoB8E0gMFpIeK4PQ1/ALnO3Vghnbf8e
t/iADTGxJwPrGivawmv8wQYIrmDwhbaVDNOvwVeQa4rgBa1R5HixNcjBB149fpVLAyJlYIMkotf4
F74bxpg33Iy0IX8gg3+vkjes7Kcy1h3gyXqbvnn9uUSZvH4VmDVi10tjVqPeGm1tHSwW/UJHn0Pe
3UcOYzXHuT9EE7YuztmE11p92UCoJeswN/fc/Fmi4tQQKMTV7U5S5IbaNKFG24puH+r85gM0TPPY
ABF/iGr2l5Spy4VBtx3KNkTjGOAbwe/ewGYFRU7ZQ0oH8Tzf8wg5VUdIIezRlNnQ+6L4k75eehd1
nZns6WrRPkPUVYWcYl84qiRFYC3am6kB5AysYIkoKiIxpH6UjdID7PYsfLNOzdkE+Go7dzKKBwv4
NA94sDpOkr6DhCFJpW8qkJKEwix0Y9wCjM8YNoGVMd8qYnyM59MNrSw8M89lbxB+xbawTBxONLn3
lT+bMu+FbNuDXiv/QakJ5TR/tKK9SKlEp0GTNuKkI5HdCf0ofpGqOGKgfJpvb0GAVHBzTVcfm3UT
lgltU3PWlTLGOhAOq32pK+m/tJrDp8QigZzXUoJgmKmvjULuCQyJAhiZaGlzyRsPT/V70B+pLWI5
WQZLcqDlwSPPpBcTUrhzHssw3BQPWaJQowpak2oxrCHJ/BY7/LeIr/k/yZzmSzleSF6NYQZrJ7jF
NJe+ySUbPBrFT2R8PU9BGWehQfXs1eMrF8ID5E4KSj7K3tWN6aZ+HedVPE8PROh+fEp4uJs6Zq2E
67OFmeyrf2i1pTVzGdK+3e5LdpJMCWwt37xucisQv1FMTV7opJK+urYTs2SbCmu4GpcKtRwdJPDe
yAvM3O63r2+FQmKAvpqIRTjtlYXKsl1WAn2Pye0SMeCWzxW7hsjbmUv8pmL/DfR1MZpUiNAjoKf+
ghwri5MJXKFEybg2E0yaGMCUEtd37/W2QOiMujGUGSoEFnGgvQCvlD5k19Sc0efPax8+qcDUGsPd
S4rKYFDYdkx5nF81MvuyjrLXhpCz7PQbtBmykFrC2RRzEgaKCiedIWsNGUCd5miFh2UOwfLnsJv8
0x0A/Y+28C24jrCDPBDi/+IsktLGSY4c54gDUyBSXF5fLxdgdKs86P4Am239sxxQK8vckA2ksTIu
YrMLx7keB+M5V3dGOcw5Dfb6bNZYj4ilYJZNP0GE5zD2K4Ak0sZUvI5R+Q6mmRBDoklb7yFArKhf
YlKPjDuEu8NH+aSu7Cf/HNoYcjzRDw+Mzt4qW9aLMtyXGfkGlFo0/Q9ru61WKLqMfpj0c52vU3bs
twLYQzJ1sFiWYoh+WwNuM3fDOdO/eTy60RHMDX82nCLwlQmCObU66qzp/Em1X5VZRjEaRRTsI4nw
t1F4NeyvgfvZuEbZzzIX6RIBis/+1JtO7+wdrinWh0eclSONfrRworvjtvqvEVfnRebQ+W0ZamMJ
wh1w6cd+xXH4yHkBsbUCl60dif84o3gZTAfoo2vn5lAfPpLMDk/LGA0/qZbguwLMZUAQf5E+XQ7O
9POLfSieSqKpAhl85I0byCx6b05WK4SV8BJaFSLIlzDtgkS8jSMmnwVhXjzUQqjl4u7K2alccX0w
HV5L2dSa23FRuETSCo4fjx+3iMqWliLG8Xl+zHZWsnF4tcnsqVUuwLNvE9TSAKvJPHN5E7hr7H4k
mwj6WhITUHadNrEjnxoj+0Rr0LoYCi8mVf4eZuFqR94aD/4JbYVxTwfpY0FvGZd+zBjfdGk6Tj7H
AsrmVnP5UjaIYdptJ6APgIKFhtQjEenodTkfYfXE7weQo1mqHMt7akNqpc+ORm5TxHQKDdAkjEcI
fksj3OUh1+T6JjBZ7KKE0W/QCX8d5oSmL+aMV4aJt2RIgoQAQNkgZfJOzQsglOYbhEYIsGDkh9Ym
vyp2bOPaliU2c42DIRVY8YGzXdfqOvf8OUhOQQMAfBxk0rXcxDe7ZsH6aSIDhPZNVJUYp3p93qHK
ZDYqX0/nRkwcmpiN2s3wDDbl2kIMjrMhIVgZmV9EVgI16HT5dgcAI7CxgCL7PSwfMYwuOKZ9P276
MSs/WTVfRzGcz2xeN7WFrJ2qbfFDOKRmJji6B3tVj17Her+UXEvUnK5pIamtBlXWYxJWFisOvWZ/
bqOLVCIQFJ/EYHSO592tKpORF4R/kRFeNtsrQlhGyWCbfVNyBskl9Ggc50bVH2OK+mU/WbkbWmaA
xx+c/mxwbN3hclXlCrzbXHNvMj3Y+pa9G1ZNNGOFhWlTC3qqoTK+1Bziir2iGpWBCjxqjY/F9Jog
kzIttdPzpReZa4USYJbCQ3GX4eefrtVWdMNELFPj51YN2UNRoabh2pXB5IkaEahTi4yTcoLhO58f
tImXaC9KUDeuPMnUQ4VG5sWH+KnAaIgd5oWlxJ7GEvgYyNf672FIfEPhF9nVFOl4n0poOBRDBw5k
nOOJns0Cx7fEj/EGePej7OH+K8+q1W03AEA9k4pxToNbZ/9uB7PHfMcg8YBeJ3FyEg6S2KCy6618
KYOLmaGdrvyfLAwU1AIeGOZbuB9kva39qLdQcFphFMjJxgiyvqvoNq0sR4lmaQ3VsVgmxd/3B2Zg
/yqK1hJQezcKAzkECytqFVKWqdWZieyWttqWMFsKAGu/23bPZwUbaK4fI4cy6GhxP59igudhVPGD
jtYhwWY7vxY+xP+8Ob5CrWbiDXhvEX06FxOEPUy3DEAja5ezu0+3wHVb/I8h6EFa/aXRBQO1ZHGj
8tXV4DxK2DMMPSutilKVOjBz0+WPnkyUxKBOdlga8NZpEo1O2G26mOEkNYkYOrlCgnS1EqhkXHXZ
uG7++IeB97nqT96U24aJlIFmAi7mmjTaJ2GACWt1LRyXCTuhIHwVdtD9m0L1c4Sos1wkENikErvG
91uvHYHB+xfz6SShsUTDupVBN0P0kXD0er6s44imjYqbKUVOGVeW5EGEFaCTZbohgK9C0gzq8Yy0
7qp9LRI/I6EMVkIzzDmhfOKDD/Uyr3uS6Lm5kBi8giqL4ENNz+65KBRKar+Q0HSr7gfG/VGQwoAt
JQqzv4kJ91Kh5Q3khbvlkaqKZ0JG4Vm8MKYyZKTDxcHkzDwXzS1hNnhARrfFjCLQooCsHyefw2bP
uuP7MiSzvB0isTGEBdMb0vO+Vm/0vmm2wRVJ8Fnv4AOVBbxa6l7+rmx79BsK72IxAe+0hA0ae8Il
gleyNOzrDDXWlmOCdfxUABZ9UZfBAtFumiaJ1pJZz3r7anrKfHZ8xsUY4UtZwxO2Ssq1jFgCly+s
HY2cLxqAgHqSTaG9VYAKVJn0T38bpQSSP/0nVwXruoz6pwSDh4HIT1eEjyaxguXpI7qJpUUY4H+u
4DVLgXUzU4lns3Vy9IHgHupEeXR8WAGpGrfRt1XSiyDsGOxnEJXxqgDNj9+CnBXIW8I/Hnn/UeG3
99nbbP5XH5J5KP1oL3K8w17Kd0AnFoimey8AJJo+ZMm+R9tKZA49dKa1AH9jNBojsG1dGmlVJ5Dt
MIIhL2cxA5eKwVLn1Mbl0LhDZU6IimgmaeJnAHdQqR6Bikvfc7+hh8ONvU5i7CgIpeCrDeudFtsr
/OSzoI84J/opEjsQLpju7i21BAcTbeeMKy+V/Wb0TU8KxGE81M6prQOWGCzcD/Gv/eDWywcnVZ2i
YySinRiIvRfG7sO1uHfRQzqS0F4YnqkYh72VZbh+BxUAhcWwGYL5Her3BzMF8kKthgrrFUl/sKGU
UPO16gjzZNJRRC5xnAWYuFiuWdTJ25geb1J6l02NFGvAbUs38rQQj5TDsCQ0zYD7pRuwcEhiukrE
ZAupRW6PmL8BD6uLVWv+RheI2flJRlErMzbF1PPD3miMV0/4Tc5LlCk7aAwYqLn424bdxxcTzvVM
e/1dSjFAHvgZ41Xefjx5aH4AXFuEx9mOpuyYQZ02y60Ab0mS4aOA6SuRTrGXf0ZEIhrcFxLoTb3U
buoD5MRWrvciS1XcPnDE5zMF3zrBjd1u1lwgD3iALTC8X8e2wlkZxr2+HGTk0QSUM5XW2WfPbZ+W
o7xrmkQg2+GV+9972wAX8a3mpeBF+kl58Tw/ny3OXBeEfBTF8belSxDIIbrdCIUkJwd+2w4T+g3w
EAVzerGTcxIxbnuOudPiHSChu00KS+XEJopL01AOp4G3c6p4LKkpdQ2T3nGXmS/wO+8qGMBxa98n
NDfk/rMVw2tWm3CoPVSCbJI4aDeDdzLpvDGm7wAmk/2AEgLqPQwfl0Z/WAxdh2eWeizohYQlv924
aVP9jRSz0Zl7x6BQ4pZFTSVlC5ih9MlRa6b1CUEloKf7mXc1iTJ1x8kTfGUZvjnkOYON8FkOOt0W
sHi6Clldy8BDXJ6QETGj1RzKVzJmL9c2aO2SV2RnURkymGrDQ4fdFahA7XLzhMlIoPceAWhZTo6I
lJMydTJkG6yCeEPglC4pVWTuNSZkUK4MsH1QGfbKs4RiiPpc6Tvo1ZDnWqBgC6fWpI/4JDQli3Qp
wctuo+UFZfcwT0GD1bvAfd5sMEIBV3k5EtbifmAO8zqDo4AADlXbaCMUK5kpg7Td48jPTyZx+Iy5
0lyQ/Dj4U2ioKMBqhr2Frst8PErv6kfLg7dEefcbsN8VHr89ce5K8aXZ2pKFDOhs9cGoOcG4bD9l
i8RjUBPsSC955J69Vq3iGJilNaWKWkueXByCvgmrO01nm3WRFRXUYTIfix+zEIFI8xEm84j/uv7A
it6yOmmoi67qSF9XxSLC4MXl8Cd6jV+8hOCRX2e6v1OOw14YD21Y76sAM6SMW4WBfrWM/2Mib/fn
4NC2GyjlhRlTrtLvh1U0hW5J1/IyXvfAHFUi+dg8nmuwGNUVUznvMFxQUbEYYZymq95uxYvkP5hH
O/otd+2gFNJuZHEiXWfkhC2qt3uSX85yu53bhzuThFAbihOP2pA1Hj6T2bNT2g/o23+lsIVmnTqB
UJE1uZXf+MtkrF4eB0Fu9M3Ua8xXX1p3TBpTOJdgkJd9iSQ+88nuDOV8r82/dIW7tiTfZBfaqpV7
29hH6VxMydShA1H9z4JTL5NERdAOPk8iUy2G1Lkv8mLkJ9kcCo6BJoKIIfsPRgwG8i9Ww59niwTF
g+R+JVA1b2Cn1gWbdEDrEyPFhN5prCqSs/DtiQxXCS0knsIxr+yRTc34DGJCRF8Vm9SRtynR3cbl
4PR1bmsCDRyfzxr8bybWKYCABRN7SKJ7bnYKhkuFm8lX6biTaAh2eXQULM/CCC1aUW4/XrWsVidI
x6wKMbrJE91yE3EbkOtCYQrqAfv6np3FNUVt/r+1v+8Dl5fBaLjRqix/QGos+AN3ajTxCEmPq9Hj
tRjzRSXQeq87yQSwgZK2IdFtMBLOoX3rqV8j5Qf+jLN/T+AnSLNpahdMyqz/q2fKuRLCUs+ENKrK
oNt2VGClQbFk19typEWIfAglnq9tBwDi3zi8nzqULP/MTjj3XGcSh/Kw1hpwrI884i2nk3xG9nPh
59yqUb7CK9qsKlJSuj4mEFySRRuWNu/WXqq6fuZFWydW56I/rP2mZXBCmUzAcgDBeyzF4+VlMcwB
9uTRKZ4e1ZP0dcWind6Bhw1Gl/8hsE2lFqZcgJq9h99dzx/a5z9L45K8MX8Y3b0orOXm+Bc6F2VM
Uuu74n8o3gOpJ0oyZekcL5lOf1RSnI7nERHB9zqbQjhR+FJtqdrDRkWK5HFMwJ59ty4H6fRgmJI7
RWEeVpa/v1dofDY+zQlWpWihUkAXA07H9ViG9nm3bx20Gl1ESQueOKpGj6Kyok+wgPCKu48I2Lkh
9eXTB4+YdIKBHoWXoUirTrHWTBgXnE7EUiD0QgPeacGfhbGvrvgNqS3y6Abz/xZ6lh3KvS/M6oQt
1VHcCb4N2sAPJUVrsJckAdbsxZJT2LIUkUe5ye3wR2CGnGsJpTpMIzOcq4ptkpOp0y/vj7jKOrK3
x96QnkC08mnXNkAUl5V9Jc2KGBPM6joX+CbIR7zqwaBNXb6ORh0tS9WbdQHsYGdJFpmZgjDJBtlN
q8HZtuN3BDCI2OMlEiv7dTv+6mk4TKR48OMRDmUya6ZxtwWmno5ZSiJSKYwWWv6yTYe/F7pSyAaU
VIeptFX1LmJ/wM7kxVleh2YZTVFPvL0FNwlire98YyRise3voM5VvQNuD7b9JQ1ZPWB1706YESOM
/+L04bUurf4r7KRR2H7eI2o/Zm2JntvZEefBD99fXO+886N9lGFw2EFUfKBpnCd4e5VvkoKJGAqJ
B8zBR/hPpF6FZByrAgh0/UgPmjRZewoQMs4lGOr7DJs/YI8vKocwv+VuUM3Rr296dFPANNRgWhru
l+kdOud+ofNPpd7stQKzTfDFOlTP53/Bu66c4dQ81Tr6sVlMkDH1nuJyMK7COboib8qYXhXDAd25
DihkNa3wJAmvfnhWzYP4OeCB22JXrjXIjbs5M5qV/V3gbMLRCrN+8VRAp9+tExYc3psT49fwctuB
4FOfVWdG+ut36yKz6S9NYX4UCWhnNpS/sBWa7H0Hw8OyXzGClrb3+fWs9Oz5gnvrcxTXlOEgYTR6
uau8phNlc+CLsdq/EtXCvPfkSRLegyK+7HQUIK3MvyGC8I1+8cpJ6xELgFfiNtFjoUlCHQ1HasYB
UEJUk13YErEOK1G1WZFYgtN83nrpYdwbOajIouUM6sXA90iEy6sH4uzPBECJH4Wa5DwHN7FrcXwZ
EgDjx/fYaFgaDIjjB2e37m2uBn9qA5zn7LnWNuqn3lrcBDQf4CUGCD92NAh4hOKc3n+VEOcICWFi
1YJtt4gL/JJF8tQ2nNeZEjYEvBLBcQkKrMYG+ifZ5NRHA/Arpo+8gaXIWHJylpJmnHiVX5nYcaP/
HROQMxco6NNq5dPrFYPgqeu/Vdx+PFH9X01HKvCka8KmW671Yr13RpTOMcLNKIut2G/EIEWJYJCY
dx+MsVM207RBRO5hl49lhziPl4+2y/PppY0GC9hl4OZgvZraLLgluIHpk7Yc52mPW4oyFmsOkSqH
mZV4Dozqcwj5R6NB9oiy5M0z+oCqkv1nTQh4hkYlEjKAajHNpBmwvncvaxh9438Fkhj1wvs4hJQO
DaLJ20xmEqGfeOLmQtI/Ap9GL1bqourjOfsuAah5CG08dY4Bn+R+zsvq1nWVKsClrZ80TJnTX9rR
aacoDoq+XtyLDqbBhJ7AZJY3NxCL7ovtMZ2g3FGyX4/xm3PSvtVlbt6VaoGaap6nBF5Am7EfxSNA
yyogDFHwNUjXGLc1m3A984UTaxpGz+MS4Yea1vzRIbqvUgg9t/sbu21MuWilpKlZEYB32JFna6a7
fms+neXUgtHdfj7t+BOKKcmb39V+9qHzm5NdJ4l1Efu14LGFYDpvlQ+HRYbhb86E/w1I+qWrKlz5
HJtxi7z/XlB+27IY2upaiNdcNLZJ/fUBr/hvaLHNS6erZTLyI5kUP/ZxDT9+cTP0qsGpXxhqJ19r
R/p/512J7LYkpcoZQzAMEBTAQhzksME6e0d/FamjCHun4H53/0IGEJhZX2w+kfBvBI7zlAp5LbFo
utr7Uf1JZAPh2irLt9RWDThRuANmF9xcAOh56K9jMdFDKzhpNsHjQB5RBE3L4lbbQN4wELEe9bwi
xcBLhSwjswOVm/fOwXspDHbSFoN4j5UWfuy3B9baS+QidTdlsWEL6BeXFG+nBTCP9675WJAWaST1
C/ECzrbOuOBTvxTJKWC+L9F5MdDdBnzuqmPNV7skwftsh3E3Ozq7Dbb9M3hgHzPYKN2EBoDMKDS5
pLz9V62hFVjUTExayd44OYOkSTbb50IW2V2+4gxH/8mpkLg8xsISSS7jHdg/f/SMkr8U8KrjW41q
iSws8a/b9S++rHlBacCD9/WqxD9/dYNQnin61lgOM4pCzG/5uwB5GUqentHuYZbAK20aZ1fVoG/H
hevKephGkIYPMWtXp8sjzsLKLDtEZoSx/NT60cmZKRm9t8vlLo6e1cKo9dBVSu36hhMU8tnRKfnb
cwby4SOXWGRMGPUZkPBaZPaAx9NyWQ5g/UdwDSEDE3wsPb3hUAzx/IpSeoPlHtaiOz8dEnEDl9WW
IP89nBvw99SJqyb0fTmgi6TprEs2vruILzVfHZWEzitf0QJ/tfEL/Yhi/xE+m/XdQ075ERTVEVsT
NDeANF6g6dWlMfwtuKbOidfRrdcRaUAbj5eXV/a3piKlcSKdT3fmMesMEtOMtPECj1YxSpHjtElS
X9IjCwiWBmw5SsPlPYBokgTzfzhMN3eNMavTmgZsdyZzClblKisyvsu2CRipvBJAlQRYl5NUEDJl
lzC0ycCq3uNSQuo9JvFCLIwr/EgwQ7d4gbaFL4SRbhLkG/rMpg1G5HbeIJY+UlxeECjkYNy4WtM/
12r/93qeF52OCYkg++Q92v7aAQO3wdPw8JPFiff0V3c0ivMQvtCPdLO2QB/W+Cczk+HQVb4wiN7O
yjVVUwcKxxw+ox3rzmy1eITphieY0oU2nRN6mzEkTZpvhzTVdl/D0ZSI70A5UoaEqi0a5Uc/h2jM
B66qgmsafuLaPR9Gi5jbbIkmadvuqrs8TkN2jE9mfkgBb+S8QS0WzXVbOMhHS1Fvo53GDbsZbfQs
EUNkJxwmBM5CWRiAB9xhXKOUTvJZCN4K9ohFGZjbRRfrbK6qzPegBTFQ5Wwyv+DGFiVLsZUZFM5F
yTgKlV4mdAso/ydLWf26VktUHnMyXNBL6mtI6fvzg48dvlXMYnqLAEze2ysbbgy+TExf+81ZSmCR
FMqKyHcUNvkOmP3HkG9zds6I8H+lVB93gRMD6IZm/RDJzXf7D1AXvu7tUAux8/We5ijjLHA7Q8VQ
LHEyPE2mcxo3AJlHz4icbRJpDHgzVGRAQhCkqhkTF9i8MWb1k+2Rr03RjM4k4lMeiWvBcTI7eFui
9M1F+0+94Z2zRH98IRaXNhhaQTvuP/Lq2IM1si5Ig5MvXUXqXnPH1lU7RFaoUs6HziUgijR1M291
/2B432Mn9pOXWpfaNtTE+d6zOBub8Flo3Ec7dofCWhxfZpJJpu1JOIUcuYIvKajGvhRN4OipYXNj
n51LNBZQQh+sXUfakzVw2kNEeZyMnJSWeY3HNkq58NvKze7SZprPjFdwLxDyCWoBQe0DV2bPahFo
+XuSTvhclabjUDotrzsvGYVhWQ5VijJcyZLJs0FTqbvnTzv2P40veSpmi3zB45fZcbadDQ4v+P7p
dSAw8/eGgNPJnhC+6v+LwWXuRD9CDTSddtV8pVpwug24VICyaYhTSdR45rNM1Gkew8HvN8FLUSuv
EOxOQIkX2F79IbfXZ5Qfjwy39tbM2PcvH3iNaj92XQ87xySen98a7C6nOokdJQDqX2Ic2+83mqUC
Ych/XX3CVafQ8IJgeXtSvaDsvr7HFqe+Ke6gx9o5d4LU8n3pxomo6IuOpYsaMajsrfKRsHH8LU96
3vs/YfBlwThY+6u/XXtrps+urQaU5jxKzH+mYit7wb6lVzuAYjMGpKbI957QXN0P6SJ6i2tWOt4N
i3Hi+4W21qP6D0DJibfUmcoSxQnnJNAhCNgYiHHXAwNSW/Kz7wWl5RdkVfmr00mrNXZKaY0tjU/0
uYoGM4jTNQw5jqadoMWPQKvt43r1xQLlCzleAUaqGeCA0ffpYFWQGg/C03f4t5Vl3bYbpOP0geg/
66QbKrq6NZW6QwEZurYX6U2tF6SSysuPD+y3Kg+SG6brDleKSAG1RHXgbcnhMKhikg5CD66uhDB0
tTUfCNKjJ0+qwqf65wGNAmIis3IUSnic/hvJVvaiL49iGz4v7WeWXogV8zHK+Tmz2ZjAeSs+PoYY
AkUY32rGkFKsKb3NTmhP++s3ykXw9ucXzjd65pfE//lHzESC5GUJ156Q5zJM4Jx09VlAgk6qm3Dh
W8XRJ3vhRn9mCUXcJMOvqCaVPvrrt7Q+RPX+X1lInfJHoyox3nIJq4d5r/DC6PtvjQQCkK9GkyA+
fe+xs/pTnlaJjzX8sOvDc1PHodO+JgesGqhMgf9/nfoDJMzyxmzTxSkX2FPRZKaMR69eyGkuVVSg
QBV3G87IGAzcwv53WlFE1/bPLNUhDFrYt7qmfqYvaBOCObqzV6TIYcX/9S+4BfZoLwcAVyugXrtC
9BhTsS6XBofTnqRH9KCpCyeDR6geiVoH2nCbWn6i3nTQEhgRLYcZjVIV5QHkrEYllIF5jLLIulsA
5Wzk2psX3Pr0DBHV2pzti7PLim2wHL6/QEKHUEdu0qS6mumECa3LTntLah3xk/FBdpjNfPPWTOB7
5sqejbBRV5kJDEaUGj/9+fqwF6tnQmStPdfmS6NkZZpRiCr7E9RFCueT3n2+mddcLEZVwOqhvIoX
w+M4ScPcOqExmeMakqYkog0Xz0rl2g3aixPSk4puUDe6qZJGgIxUWcv3zLh24z5LCQLIrxu8xGbn
91qMWQT7kyAGXd0/E5/MGvT2GAteOJpHmeGa/K60Xmv9hNNxna/YtEHqpKjFfrfsmGwox8bSBh8V
oc8iXAVzZcexT6qef4LjJVoGeuaXFdwDYevqOyDMFop6l/O6kvAtlEt40t+Y7YWmGLU4bfzSEo6P
IWZeuQdTAB/L4J0eq1LsdjzOiY0tiIxC+j77J8pxs5bmCAiRhTwJTz5jkdmERRRctoq8NYSbUMKJ
eBMU9vPvWg88iQOk5kN6OnK4bYa60vzDCN3MRZfZVPl/6hxiGmq8SW/tv3903Kk1WslBAEhhi90h
o2kgmNX502DMu2x676JZEl2AThjsxwLVc2ARg6IUn/453RoqleV6sGGb3zGvtci84dZJa8pqXu8C
v44OcUbCCPJrw74FOQe+qfeHT1bVc+fVrJv1fmW60Nf0+3nhN9T8frRXP7HOHPX8gPkXe4hmdGB+
YS7AgCeYvYzwg3ARq3VJSdvD/3/D80kZKw1xxMmr/GsEnRDvBZqgP5/44jueRjC2/P4Oz1CysYPT
RiwJ1cuz0DrDu6CZdNGQpxnVr7h1a258DcvK/fxkE43UljmJ78CKMmQ3F5JnsKBaDbqfO8IW7c9y
H9oojeOo3pub+BPDrg99xW+JDEm/t8AUX7aoVCp948bQxDoVhL2CagYU9XMXPEzJaiHtfG/04X5k
Y5x8upod3O9MlNrh/gHnab0g6aLUD/BZ+PL8DJAmskyBYD6h2WAqGOOLtG/qRzlOQtcN7IUc7Jki
I+Xx+P76fiS4W9XAhESFknyFIM0VJRjeCX7An5Wk7TFmNEEpKFzC8OUmtY77C057kK1OySgmQB4p
+D+p4uj0Hx04JNxTbbX/OKVujjVuzrSLt6K5xD9nftroc1gzlQdWqvI1d/qKi7wjFa2b8hn2xCUZ
HElFlFOHfJNEh09iUkMZ3BCnFgzHj6d8m2TmaCVBGJOmsg9bwPTBpaEy9GqwbIzxSq+nQFhxedzm
3ai2STG89cldDb9hkfdW9jz9mpN+FndpWEcjpj7+Rpd4bwcTB61j/TtJEFGukS+HTWx5jFfya+PS
iDU0D5AjezotVRs2WgEQ7rH90ZiwqipIibF7Ohpyg/I5RvWDLEJJShN2JWbO59Z5YIoBh9c0y/pR
yTzN168UtpdU3FpW4OTk6DgkFOKAPDXKbWJbPlMr0tFFmERwWq4/jSBuSirmPvovGwK8v+B6ifss
Kt/0R8gfiwF1mT6vd3kseJ9VNJmtNPT9MmP77n/2IsXbunDTu9QWSY4CZnD7eCSL38mWiQISwlMI
KvZrm/ndxBw/YVUIGrIpF9dZHw5g7cMVbA0qRi//RrOGZ+/xpnd9gTpt5LOOoPt0428A/ixW1n5X
NKr0ozVlhx0jx3MbN+v0olK72vZpGOcJp5k2ZDVADUzu6269cdGyzthLYGHpORZJlumijKg76c1t
zCsjbc/5AsPdqKZ916cTuvbHYAloU5aBG4I35G/F3BbGt3XyOT2DY6Ya9QVJO57y05zMY3mwCFcS
67TKA0aznEn4RU7TdpabKXHPUE7SrriFVEKhrpI8c73NbJ+QuTyeRNJK+EQIT0NkkvomTnJ8xres
fWmYARAszLB4l+4P3/zrBN5+bLnBX2fI5r2u84Dwt52stFrTro1P65k5bdMPObGfNpAjbq6u4L+R
j3L783vvBmlTxvWUXqGD+f8+L5EMEtGOoTCwdwvCNAGmY1qU8CU8cO42LDNBCdoJD1S8Dt9q6qPn
/McLmLp+GOBriAYxGCi4DqdPR/YpQm9TjX2adpuBUO+OZ3m7djgL5Mb9E0UyPWvIQjS6xj4gfjNd
caGjlFGDbDuzUBf5HKg6NMzB7HJeOzgbTLGNR036CHfJfDJzro9SxgXOMgKIf+ZAq+C6R2P1o5ya
xC0j34KQ8C0FUeN0FaLhRULdvR/gfOSaOTf5OnhTHgbCn5Sd0MIIYtmhysvCz5Fi8Mwv6Hr7xCbD
6sCuuzWr2nJh0/3YTqg4015oFgBSOkha32va8mFy8CzR3eazgYU2cvbG7Sz6rsn2LYFhsjaf5UpI
y5xwPxItbMY35v/eanSQ1KBinu2zZJatHgpM4Ggf+q4YpCMp5dTZLRFoTAzBzR6IoiLaN3Lgm/DV
w1yPSLmrw973oabTRInDQ7rAOHMYASVMgSRVTNrZKFVR+m6rVstut09GyirUmprYUqQq7eVMOlNc
OpLJYYdMrBZGUl6q8Pp2k5KzdZE9wUtnKL+hpfJd2/ymIheFQS4/2NQ6TCcaPWD1ZWxVvIpwiRwp
O5R9wYEcRiDHy36WBBeUJ7by/FJDptKz4m6cLqs0RnEjlgoIKNhmlf3aZ3tZYT0Qmv2Fd/lomZMx
+QaGITwIIMgyIaVPe6UHDYPAqC0servlj1eBysgimLQuDXxuQfw9EWh7tAWvH6OK0NdyVwfgLkii
PLuPJZeWGQdYhgpxbXvwLaadA22MdLH82tH5ZZmq5xEn10j9M7io7Q4RcfDlH6V8YQwsWF11cSks
GeCWJ5Vu4LtLW9ieP0srd9/BZ1KMj+89zOe65W5tn42LExG4goCjJanhynzJ/on1Wyz2hRTY4qL7
iZmV9SaX1rgSLQNyA5o8pbPfpZYpY1M7OpBvQ2EDAaOIQ5EgaXfwOPuJvhN4APGgNdp53QrqeyGk
Bvidf6YPPdzEodslikpVwY4NfQiXxv02p86/4ixZ1Pdmz9+bCqcl0himOMZk9vaOb5hXwgPUdEOl
jGjSpjCM/kQ4ZbFpphPXbwzrcCcj68zYSyknuy6gPpvbY7tdZM6//S0S9RfGKRApaVYFHIrewuSN
6NkRn8SktdQRNXGdSiDB2z2zNbWInSbzllgJ1KO8Fj4E+VqxqBBQdPfxd2ulriZtSQm1QSzKjfzI
UWuXpfOhLpBMN14x2c/ieUyIaoa6sMx/6x3w4yPe5IZy6D5oCknNDIC7GhKnf4BgVdIZT+si7bIW
28vKDGcLQKYsos5gOy3LrG/1IlPfAJBiXuFKACgqq7ZNFgk5OxPmabm+VX5Ay/Zaa7gPtIzrBFyK
cCEKyZRZnTw7Qqr/CNhIgylaCnpCoUOb1s6YtkY4XiGfNtdd2tLha4MLO2Sj3gpJnnL15q3w+Vb6
lEKqNcb8JgSaAdO16VsUHtiW79rrkxIvyH0JVZQ1YFyfOu6H1VcImYHuzV4NjDwlim7p5WsfIG0k
da8nIzDzwiiKB9t1FJT0KwGOxiDN3ORxH/fdPM2Ul31CvXzZ9cx55rg29OaftG71Kb39GYa/E7lx
uWv5zEdW7GTP7saiWquZ0DHiKxzQFtNsMAAFW89dyzQM9xqxDrJPiGdW0SvvN0ssKVkMw1xnYu6o
1J/YsUwC2kO8Q87aWYEVy4qippadB5OOpT6i+ZdFoxhQWDvnnSrBGhiP3i8s5RiD0w09gQTzGm96
6m6CIxlhGZBqcCOrC2r8apSz/uwfMj7cPMqdiRBb3iyi0gFcGCCablYYgPHyNqPEVcQ1WLQNet4R
DAoEGt3KraSoUhW5wSCzoUzzaUTrMxFXKPN777mfmqqf/uZuA++4JcyN1w6qpsRZfGCvO9QwGBwG
S+C5yTW2SmA7DYoaGVKSGvuq+lqXIwZy6mX/lG6vpXtXCgtxCqvYErx4f21yyIdakhAHM9Z7yCyt
nV3umlKkLVv46IUYrgS8E3+BxjSh2QfIhRuACVY8ee7BgkdROUu2R/gFNeKFI9J5N6d/2G5mFibe
vQsKU8HpbtnGLB8HbqbhR4qPZSDDJhk6Cl+O3Q/0O7uogonTIYcPKq7YSJFO3BEMiHOzFwKHHwfp
JkhYwBF5F5JtPBr3Dx+lHh4qsuhJ0Cc1Vcr2OtcL2P4mb4ZtXeHwqnz2MlB9kqNHtsJs1SbMHX38
8/MVeU8QOU2XTJV9RXyBB3khcLzjq5MbMb8i+1EgVPj6f8GcmQKNw7ziiqWlx/ygfuR8wB42F1CR
rWemt0ZSPRKPXsnDHYW9olMzeKlZ73Vh/tufSckat4/uaLQ3LLrci7ATNYb1mcVB+Vd4l2oRqV2X
ksfUbRj4sYyTprzA22XpivgDBYh6Kh8Hc4bT8ip3YUrRbOUfmxAQZlj0ayibRJSIdl/P22uI5DSp
6ETDmzsFAFzLHGKYWCtYSUIR9i/zS7dgF6jsn5n5sHESDneuizDUBAwD6Klyo/a52PxviyTu8sq1
fcx157bqsVIc63eTob9474EFLJdF9ZRgR/SL01g3ztYDwbJDNSNEh8nLqAbHfRqh0ErR26ZJBG6U
1tICSzIukBS0sWNsK9X9QImz+ObsEmkfnvBYxGBrooNe+G3DSmxiQwx1zULsdrqJ/+0qQHUiSQ02
p7BShf+8MpfVPFj1j8zSgVNJdCK8ed7xFoE0/T9SO8z/Cu+L9zEV4YeJx0gxooWq4hhrzEQcMMam
SRwgGvW2ysKFfwmU634fx6Y7Imx7svL+oAlhbp8rtUJcBdql/FOGd4AC6rA89jTG9gFdjVtrNffc
HEt+2OP0P3pv2ukxwpt2WKmJY74XRNiA1xjfnST0gM1fgk7rDtPaD3WrMJRpAeYlG+KfUqVhI0jp
1HrF+5E5/CQNxXz1LXrmxkdfdmQjCgnkE8IpFzFENshT06MoD0So2B0BGhe715iYE1lUl+E9w4ZB
a+/zugzrR63gu6d/tiQT8irJNyRO84L6NeXhcylEp7GkzH5BuBuzWVdrWrINZ1P7J4oFxkVdTcuI
PLoNNTzg1ubF4Vk+J31BCo75V69A8qQz/lYyYMeswEHXJ3i2hhbxlJK0fG8QvnIuyWJ5dQTFcKiV
rszWWi/k8Z7DlgAfx7it8an4IHjpKRJfxZ9+mj1eOWAItcvcUG9zpI8fLufaDey62YGrg1jhoaC2
bkxmCKeBbYgQBVCEn/2XQVtPkopxLXrEHPEkyiGA9TIlyaH+uAbpuL9UCiCNNXJ2RVgJDEpbOgIh
7JHeZXa36nQP+NBtkjyuNJfujlir46sN8AZbLi/SzF5izVr1oF8wyufkob8ETv1MrQmyTwJNAyhs
qi6QA2euGiZlvVt+OV1MSVknN20pWRQ4Wnudc/SC65yQLz++ugS7hGdcEOGofIEqam5RsYObpZ3P
eg0K0rfCjQeu2Tp/lJCjG/rAHxuACAaXAVCNw1mtqk2xjy2awAB6kLDPVvemZkAujr5zLJe1ac3d
u5RTsTsH2p0Ivybmg6DhvEeH5ZjHbH69GQmxxOm1fxSfAQDGkQJNXHs+l8bOz6uoN4i2+RDvs61M
GNKEDRklJC+TvvS+Whw3AGoQliI5wKZa//dGgF0y86ptkgCdBsYGQJXPax1Jf0AlpAsLJgSTF8Qd
ghu44nTlARbBgA+61navef0iCcmhsMv/XpLKHrJx12fCmXj5e7X46dhEJjraaSsPn45u1dx6dR4l
QAHlA1QhqDEc2oxw+V0QgJLO8qGKzjD04Fm8PIRKYArg9JNt8Dw1SEszvkCaUIBlFKHqE3lW3HkY
jmtXXhKrjgrC1mjmuARGlaksGfDRz5yZCw8sLVOsnJPL5jEtZEI9oUS95+xVUYrOEz10AlbfjwbU
9ucRvUeBZM0TPk07Pel2zkB6NolKk0J7C/JueenCybpllCuHdWGpZKtx9mSxzbbPbijBpqaw1iVI
9ImlM/8SBvp+Zy9+bF0yfHTKibwbaQ5t/Tbf+yqfCac6cCgiVJWI1pwrV3BL9oocNKIKkQF8t1Cf
lct7RiXAoDIBennbDIidC+uHtsFf15Iq4XhsRSSIc0ip/6RHyMscd/L41ccfj689sXIducXcUUVu
Kaok59zcl98kpylm1lCovrbqil321g9adrR8e9WF2R+kkCsZdoOa1YTvC8FRp4xY2QsI4neb6M5O
c2034mf3m63oynpi0E4FzHTfmcTTQMLiJgdPgz1iRNzHa9u4LhV9KBruxNbSgyazeYv+Wbq1oX2E
a2G1Duh8ZyqBUjZZjlTy4IUsBO8AQynUyd9X3pvd2P1WNc1z9MSJZ46A/+FZVRuBvc+tSEVxadOl
T9XtAeLU0Ok3jW7pKVS7q+iqe3Uw7hpNaBpbAloAhNoF6f72SmelgNsuNGunPGbyGaBSnUuHIxpC
UoQGGQFB2bOFKr1gxht+ZSmue9kfiJn89db1hAWS26yN41DfTNwFETI1uqcnP6sOm0JpNOflhqGy
XIuCo/gUeQxoC4Ivu/3Kfh9/QFJYF/wZ56/xe3BQTlMhLn1dYcp9BxuLsB3QUAvXvuTio5Jn1Otq
4cVyiYxDCPRqR6zemQM0KjIMNsu0K9l+/oDscjoF6OYADEEG5YbLOt/HR/WDf1dscltFsYVqzs5j
8DybYW5XrSS6i9Xq8WICG91xxG6S9nyFT9R8NqyMDJwAP+qVhG9HjsvKFYhChXcItbMktfb+UAVf
k18TTqty/p20MCwMQA82KPLBaeq6HLNBI60lMSSPELUVllqZ6iLVE7/zZSYYiIT2Vnuni+/0wCaa
LRcsK4YluKvE+texfJ1ThKSY6wkYUD4q0H/2llBoqt6l5t0BcY/NYIkCgmTs+lgJQiVp/psxPc2i
Qp1zTevXk8KwwmvaBqXZnZQ8rVfkYxHOlvXdH6dgvGGI42CfFUbV/OE7jUvBDOYeDBlvBDJNkqr6
GKbpxVgxzUIkthCAWqNaBElWUf0RKpn6brc2Lu54fZ8+k1REgxY9gj04yx558rB47llhhOWLTUQB
iD4pYVNt77E1bdjAQrNFElySc4CBv9tBL7KP3T0y9bZCl/nRqrqsK1eD+ChSUhTfB31bXxO7ohl/
lSrPkoaqkTG4lYx5/NHr8Qcdy5Klr4A12ixLbJvsgq2WsWBywBgrqDBiE0V03TCURbBiPvS2ztdO
/m2lGpfeX9or7JIh4os2hRmOINdp4Aoy1GH3ZcQV0QpG0u4FQRtzOH0T3MTRfs8L9X06VheKlXHH
kzV7BX4CR8EQ4gN+965nEGgELqoNV5gitO7B+i5rVhx8fRjrCpRvMuxb2rB/bthvZqGCHIBjEkmv
ByBuVvW9vWjdHuxtl3PKu+55sLlSrQl+Y0bEW65FYQMKh/jZAIDP8S1dQLgmFkirT6RpNSUGHVWY
rlrGcHtgwbwFZBkAxu9dQRkxr+CPDI4O0RWGuHwJN9CXCCvssqxj3eXvb+MKPMM9wKNQyl9y09U2
w1pbDxqiQJUVziCqVnuLw2690p5NdJRUOERfH5s46Y6z1/uoDANhAWozMgQGwDoApU5cz1CHrsaO
k4UKIIF8jUZ1q4GauS4qQbs/1KZ17CWQYcG/ydtKkZEwY4Colmb/fHgS+AXLuvQ3iikj5TkxfEK8
VSaHXL+pjN7a22bZRcAzoVbWu8Wu1MwcXGJyt/MR0t6XrfMfmdpJnZXB33HxV1syBBuHeQbh1Fkw
eaegvVbMWSAyDZwSQ2eb6bs3Lq/F0B+AiqRppJXPpVwj2HSzY8gZao2NArLwn5apLFzWM4RHPOhW
H+9tBxVYzYFFZKFBukevZauSxdnr+ZAnukNykbz4eP9VrU99R9TvtOihPzHV3zQ7dcY43ur+vrq0
WlY/Rwi8G16FbdKgDTY+4XARnu6Gky+8W3l1NzpA4Dk8Wfq/QOMDG/66SNs0sKSE982jkoI7Akm2
I81+rLOyjY3YuOhuMcgX9aDKbbgvdBFvPfbSioOxFq6J01r1qfOwR8b2SXchodoFoZCMLRt3FJBd
ts4Apc5lo/QaKaEoFOSgrMT1cjscNmCBiox5fcvr2qsYYUu5Z9DlFosJjrLwCjXtaxbG9A8erAaM
v4ZJRDLmmlrhcWVwb8EwEdDNnnyL8YaplmTOkhZ0yLmAAkmnc0XjsgsyWo3bzR68BMl0tcEs/1Z/
hFWsfllPk3ZHgQJsns4Ybq0fBHFLBDwwZEusvAt37ubKD7GGWZX6l4yxXFGh5SoB7wX/Q4O2e40x
L3fxwsMMJ4sU2w2yNk/3GKDqdDcdsSAiaUv3ggeVqSA3KIW9M5m42hVNqTqMnBvzj2LG/o84a9Or
k/rkI4BNT8lfDH8cSlB4CxpbZTtvpCnGlwN7h2w6b7oZBb49eEit+iCSoBV3m2c09Wz/8x4EsvuW
KWZfKmBJm9mqlaxFoEoHpQgmzLZo7U025RDB9akSyrUzbuJrpkLtAvJlgInqz3PCGt5A/XdeU6Dp
MMYqNTVurmVu+3DPpC87Vs7hadYOjmnF66MMSIkZaQ4F/m/cABuzbR5Kjjeolq3iuTgqFJEYCQc1
Ylo9lgV6fkxOiMTEYq7EeXfQ8IFt01/yn5VrterMRUhKqCamvVnql2oUrj81WIuB8J9eFPqJ7A3+
zS2tnm914Ys1o06KE6zA5uC/tXUhVaP3oDn6GDCgE47VjJp0fpk4XWt2mGd2gU5GDBXABh3btKga
2c2oVrxAHHB/Z4jNRIZ8TKuieLLyz2pUxpVdVHj8bkW4vaTrUW4zCcqKKY4eZR9m+jht1OJbFQUc
kDTJctV9tin18D1Hcte2FdtWGtdWnyqSJYDyuIHMoCon6yPnwXEGXpOb71DM1FFb3rqxZepfAu35
kB8ylvAV2hS037aOX5lQmGn3+CiyzSFHN0QaN71xHj2IKQc/00lanc+xxtlJH/rXprDr4H4voi9q
r7zHUXvR9pXFO/mHXKEkzTY8d3nFxDwVq3VP82T5r8XH6gNw+uitddL8qwgwB5b5+bNDjEM8ddxQ
jFn4c0dYrtLQ4a3Ftye2y8Fkg3ZJuqv8wo77na2XiJJ1MBDaw1dQy0zUi5hBuAy3ybMy47u2bkdG
cNYnaOsuGxH0WXL1TPJWoYfzHF+gmLKSeOce+WA/Q5cSWOcn1xJb8ryTY8mRDUx8Q2Zy6wokll40
C56lYm52Kx+5NgvZhMR0SjmUvUqEVxIIyDJXeLx9soElAbIXR7UTIc7/eRykskCtOnTu7tT6deeI
o6u3YNFh7iSgv6AK4Mo2B3bzhRAp1c9NyPakY+T3Bn9YZjX82NirkAWo4VQzD1j3ZkpFFk/ahbvE
EnxoQJhZ/jj603XoijMLKKP6OgLSckeXHvEt+5zcug40Mpulu1Nqhk5/DId9QRp0wLzzR0bBVXgi
4MczGcxjpiXt+CyZ9VETHT9HD4Rni3nVcjXqlRF1wzSTIGrgluwm2qGimxClnzPYvV2oulMG/BYM
2tnQ/HjmdTVHNTWKWkNmLuj4pj6DcQNewnMdRaPKneB6ld9GKCHybF3FE71W54k3R3mVxPxgjqGD
7JVBxn22SzkxPTF0e2VEiVz5lKsJ2mZDKzbubr8Ah8GSKF3fGvsO9L8xydDYhaD0EJ7qo/62P+n1
NRM2Ezwtmo//yKQq4vllf1hQe4sx/R3EeRPxCDP+UVqQ77ZPNqVsSzmDsdKoJ8PlB+1gECY0prIP
eCe59E1h9lPtbKP4Z8pK7pxql4iqOR2jAzx962bFbQYIIC9mxnnEatoHM5rGuADgo1RDNXz37WGR
KxIU1jEnARCb3+dIKNojGjT30s1xKMMUD0pLif6wmP7WrL4jsNLe6hllAfizVUHPy0O1t1rYta7c
QOevdSTv1v+UdKIyNQQ0aCe9wg5z0xt96uusLEuCIE7AU8i6Jfu2Fe+Qgb/1LZ/q+8sn33e/wB6h
MI6GDp0h0iy6YCEGZpzhlzFqVzj9qHfYGG8ZYKLkbHcO7ENf6hC1eGN4d+FDTaeekiI2Mt2yQrGu
4nAsdIXrzHEEFw04Jn676ogmA740iQRVXnRDkphjdTZFMJ9gCxPxMEiXKzANJQz5OmxTQuD8ziMG
8xlJJ8etuuD23sQ2eKMt3pwmkL3Q9WSx3XHMoFGVEjsbpIGsW/JIy6CjvBPtgU7/Uo5JSSYYl8kK
4YUCWV2rn9qQrTWEeCvm9yuoAbsJNKtG+qD446VEs6xhm3BoAgZgf3HSyzizQr+za4Rjia/G9io/
9H88ukWRxlCwarIKuBrZHSXjzLK/Sgtz98GlZn9smnTJuZuovcKYHUpHTJTNquzWQXojAddWa6zM
M1vk7ZnO8GJYIuL5Qyv4CiTXlOxyP8XKAALxxiUgnmwBsUyFkMRsyDlO8LWamZThvyOhyy1B5Nec
PffFN+SW82aJRaIAy3MwHwDCVitR59HQEv6BalZi4OvIuF/lQs+BsvF6YKbjiMwBQ+FolQWoAlge
RlchRbptZmggKjUIEmVkxdrxxmaZyzXGOQYoo0kCD+C/uTKAjSBRYGdNsvq27+U4eX+7CFUJk0yb
aPgA9ShWlV7CmyHmYJ64sWTaLqZm43hu4hQqznadeAIBmN7EiTNvO84lZNOKXW7kR2RQVAu7WDRk
5x8EXMivss/n5ROCvB45jaLSzLG+4dscKnF/cgPhCRBSF66ojSe32pnH23l18cosvuHdgXYRnnup
rntmeqE4AQAxB3fm3KBJQaPbZwxCMsfXF1qST4nyO2HqwdYrg9AqluZn/4R5+h4PwUeEJK1h3AWF
JShEhX6l+up2K5O3R3kQSOvW1EGSFNkObeBSS2RZfzJjp6SnA1WucFnwTlOwmm3tqmNZ/kdbX8v+
ntBcnArjyvRJLFNomKDXMtTQ4llhwZp7sAtMVtl6gdSlSSpUJaX4YY1dQVDONYnSqzbNRBT/M9un
fQXfAQJo6qhwRZ9RDCvD9pmVwx3blZSpejUoY/oCnbEpNE/mim9BIUY8od9iHYwkdstWcy6tg1VS
oxGj8sl6/XoQoZoBuy2H3J0nzxuppTxD4preocn50tTVIRvHiMzrflD91RyufNvulFkBIgiwMY0h
8LjA5x+XGRwy6cLKglGzYGRHgcq66Q2SuUI8nL6BCNOoTfAi3iifj3E1aRMbln2tWtIG9tN2YhQg
brFAxrzfLOkIZBKq+kKU+HOx3VFonxo92AMJnc8XiRHIDJtCYdEk93PgSiBWE33JTuGTQ5UKsknS
ghNEBJwYVOFtMONzEGxqLbVmuNmDMx15gWIuZSh8/L4uQ4VDhlb36EksRfOsyj680JVmiSKVYx/h
KCvyDo+oBYPQUCWNM7szWZCtvEypbenz3QibRz9x9ImcWRXgm+hOAXkOokgv3Iiy4Xe1qFE3elx6
AWbJ/criDy6LcRzPdnMakwvT9eAzj+BPDe//6AsB4ArzZLfh6xip3YzyagbnTqYUj2nrDKmm9qb2
RRtap/592+0WCd3vtPNxJpVJP/HCQcnKFFexJ5895N/uSHR7smTfHE0DOuRo84XFO1bC7rNvJQad
/UOwPWa5qv27YKFyFf3Konb2LA6LyWnmyPB+TR492oIziwpb1tk5YWt46ywTuvU6Pn7MfCzgCowp
0s6pjD4loDjNdpg/N9ZgZFvsAwSV8K1GqVudSTNkcpC+MuNsXsaBfkU/7lU2hWVb5+XRhheQBvJX
dQNFgKAlDCAmzmpprtGoKHqoNyGC+xDEHU4bmJanZrvsv83UPTh/QHVcMurtMD00xocAf853Xpj6
Jih8Wv4FEqO/TsLOIFndLwdSDgrB4LCaq0jgZrj4fJ+b9WUIh39O4XqoTL667M/2tQBZ2BYH3ZTV
xNKjDrfj8gUHYEO2wfL5HIF3bA1LngDm7A6Pc7w2fxTVxvjh9EatsSjIpTLwCPA8GTsp2x6uvTP1
vyRuuOO4Ow60n4qz4Rsuz/32ku4HAI/0rw4xwkj7+L54YW0L9cExJEtHkp+KSjWzH8nHzY8mR92I
EtKl3nwQrq23Dnjg+xihjFzJlH7hbjs8fXMeu9Wc67Hva1eOxh/eJ+/u9jS2nwqtDL5MYaMhjcj0
gIujAFmDxg8B0waSebfrxLYD2XUk4NJ/KRlIlo5UpLRYcGDvUliQ0DqSNNsIkqIIRVknEgadxPRX
QwxwxGn+zXuK+8ERfB44s+4xglU3R9+2jDgKy8VpYaugMFLakjygy3gvqcyalCawIm2oAAdz6nFp
8P7BO48pzGt8iK1vzicsu8bbfFeC2IBEWFBv5O7g4rF4gxEPtKvnhwCjUYP0zOAail3N0ZPZg7cn
WIf7As95DqOIuHbFsz764k+W4nQJzGl4PCBbzsRQuiJPa2Uu2Oo+lGys1tHq+ZUDv/fzzDrOzvAB
XNngvxOVrDMc+wmsfsKKoyxkZ3Gvctn1hxnq7XFlZA0CTZ+kmNa002woyy2lTE6tJx7sYVFiv2Z3
jqlDaQ3w7fSzd5gFkyh7NnRn2GNjjbPrGvvJSG9gNPdy1c+fkMmIeXjm/Y0Tc/Oi5Aku2kzclv6L
/VFjzzBkL67IWQAJDOj2NQfRCbY2SEFCyjKfwS+4LulJB8EpdTKhNS4fK7gtu2MF8TKdXvGM+S24
oLT6RcYU3f+mnMD6SwPiW39nG8xQJfiFJuIeAET4UfGuO5LX2b7iad9R4pLDn8PIf2Rn+PjkT5L6
d463WNkhsjIAUtRsxoqLnO5bjPCoISp6YEyRaigRL1DpCtg/lGv0VGVqqaxAop2lNsQ5/jdc+sFF
5Ef9dJvFdZbFNQb2ObD/HM/ttlJPN0lN2zJfhinByENd3Jd9pbLQJ7OMgF02sT3G0KkCmSkU3lN4
cZbo0N7c12nm6mDbGxwo0O5Az6D3cj5RXOcXH7Tjmg/tgsCUg/f0SXv06y1380Q8zfkfphmp3rVE
XKkmH4wVxqWxTg32NESYt3xz3wASBRYR8qMKNQCmXKPKwl0rIP/Yv3laUjnZUYS2/iD6BGsoJzqQ
spdJA28qpaP3DSHeX6YnthTbhbsTC2iWsPLzv6m+pT0FfrvzV5JjmWG7f2Zl6l2p6ZHmNuxqgmJG
vBfEGUhOkR5Fv4kkCL54zlqQOH27iMEB74hlDqFrvhYjfUJW5FdxViAFW3t+POq4EnHPuVcYauRq
sxfo0oTex0er9W8x6Rww0fznks5xDcxR327wi+1BfNMvPkv5h8Gn7gc14ttFRVZPUHlkreDvNtY8
OanIAUzTN7GmQJFderD+WzE0CaQWpKTUxkaCMV5d5r2fUCap2OqvfVl5Z2cqMTjwrGzYPbqnuBze
iptjcG7HXWCxYeMBw/ZRkxK02+BCXJr6klmEEXTc0iF2s/WCSvN0ain+OrHr6jAjuTTcH8hbFFjw
wSyQimxr/1TMMiavQDBZnFizKOU2ay2V2KAJVlDqOkBiW0dKRuw3EOzdynpqqrD/mANyTWwVlI70
m6hWHGATTLuzOneBR8BAA3Kl3HxrpLy+Dfx/iX3kxo2IecmqELwFEf5CMpa6eSTUMokCLtmABufN
LPkR/3wRBjuS8TO/nzolpxw3OUyZycnhxG6OzlvHdGtg1J36WgjXHZFQJR+a59HY6RhGNhB+WZDE
9NjJuUOg7X/weurxZ2ncnLudSohOu3T1LJDdlNQVSj9C6IZL+0uMPId696sb9fUPexCIOBDgfKuG
wzYVOBRA1poZbaMxmuVRlFJLXIeOIwaLW3JwvYWApSUwhpcvOKfAcilEKK5r1suDc41fnJdgeKIp
7e1YDiqeCehNZnDWpW0bWuRML6qRmI028VITXQ5EjwU0/YUFvn7a6tAih6fmTByUA2QOKVtxpI8V
yUbyUxHrwoVoT2GDqwEuiXthBIm+m74YT90b6ZgYHcHK70i/gbK22Rly4p0e5buAKH2YvbwM7A+s
nLp8C3JvsZpnZPJtZ9kT005v/67fdsqhXMEzsBQ6eaHD9JWT4WQHMIXq0gEbGTH580Rb2c02GCjB
KI+X7iud5Y06Cfr7WBvZCgvIrmOk8D50K3TahaueZz665qpQuUDHFF90n5HMhgFDjLKnF0VmL3GN
VTf4gcMc8bpHwqhQ0BRcmq+jt/c7Q/GW2enTrc8MXzFd8mPsY0YSMh5t2RZ8adU8FqK0dlvLBxjK
7toHGaQmnQB7fu2xLAa+qHq53Wh/WD+Y+22aklQS4vGK2gOkXqxc3ZDSvUHewCuwS4xtV4DeeD0+
o55hZfG4RC+KdMo+qBX+Mv6KY8M6Hnyzsz9veaFp1HVqy4MNLczA5SZljTYMoN8F3JhFXNTQXon5
DdDMdX8aFH+8th1W5y79VSAP506EL8PmRQpJwChr8f/RExieE9nZy6i9pDsPDfxCr1k8AhGX+bal
+wneZGTPZLW84kapCn/PGkv81UnfzofjgrHX0XkdmQRxFJF8O1yKXAC44qbphtwMOWvtaT32rrUx
ZkDo9aZMfbmBma7tRFoHve850gPZvYAnIf5vVOpJyGE17fk9sFEU/MKzjoRKSvDNwi1pF50yNkfb
KGwLPC2Crv3Hu+KTpjaNlKq3UzsGBQIMRw4FkRL9w8IDw/nukMSLvEpAlsdJMYBEvrgyAFZouMYo
z1Rnt+RJ2RCD6xaEKLZthfS83niqfkqMXSqDOkaXOA/m4T/Iegjg5Jbbcy2bv/Gp/GNxVIDBwAqE
MhnXnRLycL/vrp7xVxitMP5/h3bAJQ41ri7VnwVTbFcj+O94uxHi/7V7K2UOsZwLmaLukyrFfUfl
Y8RQuQhSfgWxkaGgyQ1d5PZoN/7UW/hiFM/v2GJSabegWEeQ6V5mHaKVEkCcglFT2BMywxgPUWBa
VBBiIhpsLY4cBA4JBZxncIl6DYLHrfniKVe7iVZWtC2LgkmY1mf2v5I4RJHJiBeGRV8064SB4hgV
9O9/HLa1b8iioQNGEaf3YuwFOBDuFOZhkmELZtCBJ7XybPdcAmZ38IH1P58AejhdmGF8qMn4GDz2
+7qug4H/0/QTjjnDPdmRZp0x0/jSB7dxri3xHAAYsfuHpTrNCniDa8XvSc+oDdo6CGduQ9E/i6a2
qmSZeoK7F2Zlnb4VwaM+1LQB7mLXczOm+YA6iNLLA9+rl13dPKyyMF8UvRadS9UKWHecXejsi0It
hwdxa4oZ/R+igXQhFkNkG8gzmFmijPj1kd7sqe1soXIKEd8cK4w4Kb7XLPBx5oknqE5pKLU/XKnk
66aPbfmhrh9Q37P0BrQxy+3WfxvGiR8HLKs02g58kk0BMHMtUINDNoQ7b/z5n4T4jXqkXCPz8n7u
L6pCGDFDHYPzlfyCXd+uS2DqVMk44n8Hac43w1LFxHBbC4Jda5OwAp5zcFp1iHb4C4JvND3MfiNH
bkUAp+nyoIXutlhMlvhM/jHAnCa9X93KKVWUfqt1w1O5IEo8gXlm/xP+Yp34NPeE8xoLcq1Ja+4o
BRv3D0jHSD0fGeUh/p7RcZcx2C5jUI9QsaLEdOy+vBdtrvCDf9cvq7QnJB1EkO5covhkYcdK2+8G
VH9xk9pPiUIK5/3djBNfwartjBoFZxoPW+2/YKjUMp0k/+V2MGy14QFEXRzRYMegiBUonunJiZLN
JsFIJWlXbW8KLpDdteP1OXJpmSH58dX9375EnTtcb6w0n/10LfzZ1mcOjmhzYrp8sA8LS4JOR+ik
4YaqTKV9RYSvbUZbxpeMG1XNzq/D5FLTs9r1E8Ia7R9YVsSgq1Hx13FMu4AOnXReIiKy3n97d7iR
5Im2SGgImfJOVJAi1iReCKWHa1876Dj4TDPKjp/xcZHBKaKsAVE7aI/bwg0SNmkJJ85MIdRm7gPE
a/aS7ypaoLV50V7xv/4qKfgAiIiJIdq9Vse4RIOD42XEQl05WWqf7mQD/7cVa4oxna1muxa+yVDM
m25R9aZt1ej7qGURaU0yaCVoKv/u9htavpHo8ftg/a+Nn0JK1z7rooZbigpdsrCnqtDaUUVaCVdc
rdpFLYx/G/gTX3xhik3xD89joenH41MCk7gV7HkGnFj8eEaO/7Ezncy8SmH4/EVLUkLzHTf7uG4k
Q8yTFdNKkHLFI3qaiiHZ2AO4sEFe7kqmNbWyJ5cuR8mg8zAmOJe/zGdIl1I0PpAYoElBeJqovgTo
VvGRQGz5REu00bOP5Snjqio4AXfkm//tJPh+UFVe2q6oEaJi/PR6ZEVOQZ/gdsjcKd4QQM3QeJJt
IpeFlJx1qIrNb8PkhpUIXFjAEenREhFfQxrcCyf6vlZoViIkMfY57BDDE/os7/UnSFA2EVe3eI0P
gukO1rc2lpQ+IhOlBslxxkyyNjnSRtZeuhhDdnG01or2Kj8jqlI6JAvNomzr8LQqoZLIc3MqZuB9
9OSs6ezS+vldPF1jbqJjvEgmMJq/vimlmvxNNwe6bG0BaUly+H5xESCRHUTXdTQEuILuABS0KbUT
5wYYU0Gyu3pghNUhMGlAckgDqwI5JkMcYdz0IDKxAUYVu7gq15r+A3FpQL0BINRey4IzGwHmMbeD
JmbbsQLH9sxck5ep7k76IYpgYxKF9HkL1au8IIuwmcrRATzDK46h1saAjQu3JLD2sb38S5bETLzr
aiv9ueU2wIIgEW05Pk9xVFUoylPw0Yw1+kQyIpaQiDdiJfijy1aAvvz30M77SZSd7I4+0A/9kKOi
zuRfY804XGxdCdgx227oBeTOyG5/hQaQZiulu0+Nm3FcxFfo/x1YfJ0bHbmQz47XKroGlQGx+pxI
yzbO5hfvfEioBjmd34krfRSZpGUBoStA4usKCwxc5w61T9jMxlStQY6TTd7Krv2493pe72R7oBUf
kzu1vU1JCUuydzZhjwhp94cVN4xsxHBHSG7qwUd2jS3NH7X19OIU0/7s1PK1O3J2PmzdZS7Gq0j7
+knXHvc36iVNDQ9fNWVfEwuxLsw7Vi3h8ML2k/28isbUmzA1GX1MzHZ8z+f9zicxcjoknp6jQKFo
oLKs54+pZnCe+kZUwYXp7BnMxMYtzPGGStvLWud0eCWflxBo3OARTniPleoZt9GBNSifekdV55jr
tyUDuJT1Uo1GrKMcLF7yKGbowu5sS03xpxJNFux6Dh+1YcIWrJOwxRs8oYf9jRYVvE5ZeeiDsegY
IYxpTGg15oq1xrEMxDaoXAgONBjFR9MmtA8bKF/RI0x0chwPW4cs5xNWVh/6fLQABlHfSoDlpqn9
ASREvzHV5hOvUYa97OnH5Yl1PTYZAO/ULhsAMJQrmHXacU9AX5Szyzn+/E6XQh8eM4DrMunnTMcJ
rGtaRctrh+2on3o2ATF+2CTU0tsK7C8KrbGLW5K/ZEnaiAK7pQGnzzIC25Q3A5nABP0V4Z0+k5Nb
ifygVKCCvoUuh9vtt+4bcluTN4YJU8sgUmjsJgIcbkaFfgYS7Y3E7sMcIMpqyKLrRiMODTE3YnaH
OTxsIUdA6B29q/SjzJl8lW74JqXHiPrEo6Lwdx23bK7s3u2WiwZ9dzArUKZPUh9n0A39jrlzY5/m
roMxLemc0jQq9KPKvFITgrL/t81Darto3kwhBTemBDU8l5vl6u9k1uHoISFKq2LkV8dUZa6F8ddw
RKMZzqWHs/5Ez5jk7TRrXIXDbEMNI3jvEZe0GzNZqeT5UggYxgAqagGsO4GyDXz0KyvintTCS8cp
POUEyJfIu2yZnnsiEhM0td7vr6iLrkrn7SKVzW9se3J3BoAONOnC9XX0pDJ6O4iuuQ2xg1YdlIsK
GkC+832LcJIfadt0rSqGWa7aW7RdzqaTJVtDOoq/oZ0QtbClc6U/Wom4Q4QNEJxfy9+IJRQBfa1Q
nQnFhCoMbnjzHPa06OphVW/lqSSp9rIcanqSEPmAvXgjU48XbNWcMO6FFw8JDVBXqOGtK3f8rYuu
hAiz+Rg/Ioh2OnYCWsAO0gC2p2kfNebd3r4NFCI6NE1VG8M0wAJHjWIu3CKR7AwR2LyeLv58Z5u9
gA8Ke8NvusYMQZNdxPPfqe1PtPwWooUih8eLJSVnjTDFAYGS4daTYcJbe6GEiFrRlSxqD4aHzLQ6
tGhoGN2I1tXU9eR2CcwNRHqOQooOL1qUOPiGucUJFDzrM7dEuYtM+njCxrnLm9VTlgCT8ZlpfgXk
nwv8vVXu18e4eqx3PBLiWvRlrnqlYl+bO05T4WO8xFHPpS5AG+dDx2u34HierEwYDSCaktmtL+Ny
e3R7pQgn7UlEfRpfWtbgXTwePOzehuEGPwA1kFguEhbP8Cvl+2HZne9QGll/FgpUXIyI4n3fNuO2
ARbOdNDJRpj4HVMB+Nz8JeCvDmhh0FK0nNpwg1idwbrEy9PKb6YWK4wLRVNgVSf/z86y0pTApiWX
18zRwmzRWFr12kpES5eHVjq0qNx9LQKM4xNQ55aSohTlfcH0JFGyzsaiZSJ2RODUQxqaNs5aQuJ6
Ymex1V0XwOdzUir22eh6+zxKK3PwwYrPn1LrVZx9xcI3yl8YFcDdXZOpKuuOuGbuiVaftn8W1L3e
qRJnzfaqMU4HEZyalwM27KDmhp615XQSr4lLysmr1N1E9VxHr8g+j66gvrXe6QYM/Np1t4aaHlmT
3Me2lbxAgu9QyywK4pKqp3zdcPfnHSvuiujU7mYmPw7kMlO00D8lpQCR402Txz0pHkF6mHXhyMhy
v79gfkx3Dqu6Kt8b0l+igVYepyiZgS1wjg7IUxReg/nt4fXTHXKCrI/N1CfnWSk3rAq6BIK3ySr3
eouxjXcbKbCTffb9Naed3uU38CWJUOD2LpEDJ0S5UdGEJXw+g6Ip5TEaQYboY7yZPv+seYJhSl/s
ILsB8xUy/+ak5iuR6Nr3KvSt8dwUdJoieGb7iCIsAiDNZ2lTALKp6y7TAffe7994aNZPMD8lCxV2
vyPLuLIS0iut70hN1QPbXkvBeAaH5G/zgGR7wVmQ8aRfZLoB0s8leJX6siQkxJngIyVi+4TiND8N
/4W78ySp50zcPUcnndd5Hd7k7E9u68PcNDxeFiskDAvNhkYKNGEbSfIDlI0daIGrISqzsAtovP5g
m4yx1v8C2kaQlsW0jloISdKjeGkIopB/Ep3opBySFtT9mkS73oTFj6QDL9+hbQgN9Xl2/wqx3kAW
ilpPV0j+pbjtK+5Cot0jzUd3uMwFQmR9YjBgUcfk0qC/M0Ep/IgCHJdcn7Ye4EaJVr24mWHQ8CB0
wjRl3upfexX6RWujuhV18fN8gX6fTw4laWTIvuJVQszLKf9oFSglIcJznNQroh9d1eOyUA6kNlFW
B08eUMpj0SQtJleOXX69OHwv4q2P03cjbSYI8r8B7WxW541JaMgQSiBDXM8rvG7mebvDbdc51ASB
vqbDEEeYHk9g5wSIPj1QN7ppmpe7GBMjdAAv+mjCvd4w/fP1PT1D0330WXEZZyCsKJryugLYukX5
/CBNSR2RDmf6E4eNW/D5RqsmI0fcIgGNtwI0CaC2Q3H2C/Cbfuh+DD+jfrZQIN/eW2L6sFVmMmrg
IJxlO3NSKXQevSYAnRxAy07gLLx3CeiRVOyf1mfNyoTheR5NasqekFhZWQC9o5wuT7k2/6v5eSpt
J5H1O+NAar2/kGS1gOwKVIZeRYgc8fJJyeX6lqDJWUkGy/nCgUZpt/SHKGo0Uu9rc6e29V5VcYoS
QllDoR5lF59lhVmd75KsKTXspd9j7fHP/vdRnPFCEo5OBqxDrT1ouNDLSO6c+Gzqdt8rEFQraqnT
p6gJPAK8v15biSaYm9vsBPdY4lt8Zel/9enlNU5l8oIO50a7dAQgl4MxHBB6pAhveu4klmJUsYXI
7IzEvgL8+5zeTSomiHu9Gy6Z4pYVa69V59n8l6h9F22oW6/e406MHO//UHmGcfiWwiNX58WoTmJH
974fslkEy169iTCbzdE+8z2AG5j1zHnu6Z9aK6d43DbIr8rAFiqTtb+X6+HClKubQAYQA5b9fVRu
PdZWXHK4pDvU+LLDd2r48tXQIqFfA/mnaRcSPVshuPhu6rejeNcdst6bKfxRkv57uQO4EJmTzYFq
hl6+85t1S4EWGvFWCGtCvMjTxdTV4OVAlWSXXYK+TlJr7kSRlBGYdzfWSgQhLer3iX7aYxUvCqc5
A+wS4J7U4KPtA8Z4nB8OF8QiCaenA2r84Rmw+8IOEE43LGbuAnWiWCq6ZAP3TAVLVTRYzCciqUqv
RbfduBE9vSxvfTuHp9nljj/pS4mzPhHd1aoiQqcH44GEUkvnAN+yw5MM576IWbncMKWXZneOKSIV
TdCFJX54cK/wZCKEgTZhGCYwQICm1U4r9jyoHnfIEom3G5OusEGVBMAD7ymZg39Y56LszXEOVOg3
Cco2LK55hHyWNQYHuXRsMmn4qtgOlLpn++pM0LxkyMV855kNNGxDnhQmlh6mWS1bVIs53exAWA3O
Pa9QpjX3cY5xJ3iIA+7wxvMlugtfINRlWjzoup4sb8nGm786DqQm2ufQGib9S0zXTijNokL8RuI1
YE/f/h5IDbSRpkfO+IcUCUkF7nGi/1LCHgomg35rv6ew8rTmGfb2rePG9S1q/QdcfELwuDYh5UDW
hZyzeqwM/UmokIVJGwJHf2S24gJt/bQEd0gG8mUWNBvfnf8hVtXNSqX8iBuT+dXuVTk312kbc82/
rQp5HmpkguSWuM9JWMa78lV0tGmolsBRdPejQRQDo8hz7/UdI/vMlvhfcV22UQRntmkl1c75BeN2
fqFalHpKsboWfbKzmXl6OcNyt+6CiXbbc+dkk6Hgh4kHCd8P0xl64QC9R5/G5ZH9sq8lL5H6nayB
ifg0fGZjmiOaiSxzQFesXM1F5Kcn/3Kp2Uuq4pVegnt6Of3vfQV6OuYnYov0syTq6arFgz+haXpF
YMYbdF0Y8BNvlw2lV9qBk0rCQmLtk+82NGWJruU1VQunh+M5VgLErml/g4WU8naPT99L48hJvTBk
vhtpu3kZkKFFWKmNan7fMAGgmKwdUPTrL++kunVzVWMXd3dLJp6JPaCFkA9yhxobwVshdppqzAZw
vXe6KtXirNO0YXnITaMR3aHtrXR6YcbwhulpR+/H1vy6AEWwKmw7dwar4XFI2fjBakP1FMx8CyjX
LOWGpj3GAPfYeuSbyw9Ne1dAnHVJDlXN8AlaRNlNTHeRA5s6eehuG8dn1GRSUorwf8qWyxG0P67n
QDm8XHEaYveXO9n+OHI329T7D/y83FQStq1/+3E80tv5c+Z/r8n18Vn9f4chcM3B3LGuBKXX6ctL
xkFlf8x+gGhmVignXYMvLkJ36RHUvP0EO+d0jmKKThGvNbZOtCyxXwrlPMoob9VJ5nBHODUwvm60
b+DhV4JvTIclun/Rs+esgEDBjpc6Skl3MlXF6kbeuVtoO4ar4nwuyNi5tuyQGKfiGz87N6kR/b3M
Tq4TqVw+lDyGnyaQSo6Xeu4mTGhx8Zh2aKDjc1M+TOeQYwePUa7xgkoBCuS/L/PbgH1cQ6L4GJPq
S3mtfUVKwiJeI1zwCqLleBp4kE/ybMNmAOqhmsNyGil2CVi18i8d4zVgwMOeQNFl25g1chKa2con
LNGC/ysn2eFDSTI2EZfXN6NRsVwfT7p/zYp409qCGRiHmeh2OC1gA2kvl2OfMktlPQ6XQBgbugQd
xdhIELzqptbR0D6wRCj3lEDDukpwy+JVEynk3XZQnodIXDlYkvXMeZ/A2NZJ8kw6v9NrGvMDR/iw
gvdQxeUQ2H8its1v6hgaPxXnzQ6rmHcRdjn7T9ZMjwP6WHA94oSTcEsljHNGf4xA+UwXXeMtlS7i
gom+48bqg0Ci5vuG3fbl1557cSAETk7HGwD/V9bWjAJdCG+rTUooKZz9jcnrTqUJKRgtyQl8d2WV
2I9zBJW2fFJzIPvpl22Ppiol559zHL8Q0heaSYhBAMcektYos110KobYBKs2qKNfS87BgkHyDgqZ
VRLNmWDiFqZ4rYi3bph0wnJjrgB/CElWxdx/3rqECEp4R/VG5qOayf7cvB6oXPTPKwMiJSs3rS8Z
TEmFD9tXTG/NyZZ446yW3EGoeA5MsGEWpkz80oIAQZhpzXfgo1Bg7WTWndxVcqJDKJGlQ8/zEIMH
/T28yNVQ8fRJ2fZBUWjx1NoxCwJ/BC27CRMpnuDQXBrCf2tdQLIVPiaLI2A7wixIQ6+HC/mRDI13
HW4ZSLSNjdye2ENl0yWpE1waj+txoTi1kh7PZNVMMyh2i3i1cAArm1Xa+hG3drPXeP2T1pbXqH6U
fkKzW6P/zW7w1DD3+3lPynhKxs6frPiJslhqGZbW3ZzM8h1c0f5H091E+5G50mlmKNbMKisWdk5h
8mT3KovgjElLPGI7qFjYQckuAFV8PvQRVcltY8M80N+GR2WWVgT6A8nLD7C6jheIvuQzwq1hUqaP
lwnYQc9GKtHid8r3Te70O7S3lVTqZUOgkpeARK8ivBuX02L8FAhWv1+CbswA+vdJAKjfUda3Sk2+
I+rzdP9fyl7DJdvWG7spWmHYveq6DGH+5pc8KLfQOuEyOxhSCft6M7xG2eQclmzBJV37aJm1xUEH
f7IbfkI9blI9BHpzBT1Ey7t9mUyt2lS/8qYjA5/QPGWIWzUAp4taliG9nAAWix5XHWTa3aVCxEO7
A/bztg+90vPeHyd2+WAes1Sgq5KsCnX3aPfL3isl4q7gMYidtuSaQ6fZ+p63pen6thkbu6rhQDMe
J7u9s9aG10k45Q3pcNTb+Mtb8evp+7Dsc70eH/YEBBWxBq+NB/jJNy19mrKYdGhiTQwK0lZVMCLO
Exv/+y64CV+njYF/f/o1IcAweTx9ohrC/+BBtFsbymOkWPH0Kc2bTbI11OvYrKpTBQD3DC6ZIj0A
QgNEipgaoDwGPSqNHDC5A1H8mXLZ1MLtBJLUgjx4AmtxPqyYe+so8IRQxgh2+6s/hFFS1yzJwjj9
J6DU5tJrYouaCGIYFCxE0DgKO+S/ea7HQi8nPedH0xfX7gaTnHebLi6627lPJLqoRO5qVx0edUUx
3UPJb90XpT929fMOIrnhnPUdqEGkPSYPxDLhvn9ip+hJBHbkkVCqbyGX1U6U5NVslh4OCGEO3CIv
PK7kkFNjOmmd8a/O/YILysBiJ9iy6WZ23NgaazK+bTdJ1Ih8jqxOc1OggR8meGfSuhJ8kKfZtLjg
r7wDkgYMc6ImhWcVIRzMGGDKJGeQcEm4pzAz7AJVEOskMMOvsgQNstvT24ZEwjD30MMebMYiJeLm
8qNpuPgKiihynJOjnoXu9oofxcnziGtXjHPCJGVzr1+m/chirh0PZUcX2miPMHiKeOPYBNThQ8AS
zYq97O41TQbpB5GTtUWUdTvO+pb+Iu8SwAn3gaN+xLUC5bLv5ze935N9lM6VJGuXlPo5TIIDJ8NJ
XgfjV3r+YHmX1xvY41+OEIKASjlXW9MLlyNmD9/lC0A9/1wgZBj0wGheqP0ZPsoNAjHu1co/aspe
z4NrNmFd5heI3ri5psMWsD0Uo+cyHYnwAK3QKMklBlEFkk4CCaLhRkZs7QdT5aC5H1D75NbDNE5p
VHgpuJGr7S18kuHfEmyRviDGJxWprOhCsTE31qm1zSXysFAHjGYgQeRFki3EVXpNo55olyNZFNxU
2P43yDHteAc6m4k4QN3NgkhxKbpEGyC9MKxI6gRBIMxfOnHeytiNvq4IR46i/G4ncs+SzOExID8M
S2Eu4UjRyFgJEi881HSwIVq2c6L4m6lssu+0HcR1YuwLraHbC0RID6GfJJBtsvk7nqoatuWyiE02
00vD3ACjgj7P70aYbZPTe8Q3985lCHdkO2fK6DG1U3MBkapHnDHss/Yi+EgsepAw7+kOYtJIfg4j
ogf49F4Q7W60buZSN6wmJ2TvwA50nih4AFkIGAUu39LOyWHfBXiKnrolYU7kFKBCWrTuUC7G9QOG
rDk1Qbzhu2B8AdnWjMGqNK60ia4BlklsA7oINX3JxnmJms2YVtIzPodmJzxVY6weOuEmgaRw9fhI
M1UXajPdihLrjFQEtW5auq1JytZ1clbwLOgvgMvqOODaEJGVjTay0uYgUs+VAXYsBDl/P2KQa2fn
S0SVdyYsY7kxiytiLF/TZrWZNZu0aVujqWNdFAtosmwLxWKrhau5aCy/xZxJWD708+0gfSD1dSvf
8Cj8TYZmMxsO3KwRk+i0bOth6H2gXzrhojCfRyGOylHx9BpwO/zMwWrjlZk4aYZtIcsYvIe6wJi3
r0uEwsuzK21/vetBF1KAKiw95XPq3n+qNii8sEBzNhuuulX+giI93QzpAeBCs8zSCu2WL7Lp4x+w
+oMpLyELHqruG/7npgAKdF8SdY/fDZj6euUsb/yOCRHIIZFmN5m47dUZkgHYQTVcj41ECdkfFVLN
44loU2bgWmd+f3CtrDKJZ/8ki9piDL7gaKZWETVaNQNrz0C/6zJ+pC/poHYdlDK/L3fS8nNLa8om
XZ+XwSkp+YiZmN9D7Au/NP5Yi03rnO2haG28VEwpVpnJomhojFKsDhw6x8STqqZt1AjUBWDvvnVK
4unqxGj3xOxVzMqXSUPRwdfDVTORESg/Vg6PK40mSpnjYbSmfZ47m7DIuQx6DGEcZ1rkV6V11WCZ
zH6Jcg+0VoIR9R742a2lacW92bQ65VZIe2fKY7CL11RcF+UKhDYXqyLbSsc3XoIR23xCMXzUuFP2
WlJm/xp3t3aYwkNn2ozc+YNXcWuABwj7vXVYy286Sot+brajgY9szDmmRyUjCTqzP6TubqSRAySx
uzQr13rftcdcRLZ8EZ+tvwG9OHphhh7vUK6fhQIHVnelOAF9+uXqKHwDP0dsrobMjnwBxKy+/2Lb
Bi5LXfJ5B4II12fk8RZpsNGxAQVQ5XqJf9MI7VbcaItPb/Q+jCDXoTME/+gmXfeAQRFUZuQRktW7
rCKmYnH+6S1ziomOfgC5kw/pN2WHpEsWG1oZj3f7ZGoLZ2T6Sk/fTktZQqv4PBDxcPcyf7gF/o8s
b/vHaaXVnAWkutkk8lPREMLibjXf8HsXUTnb2Iq7FqS3k0u44/wbYDpwIicCBWRvoySexNYnzSzk
aKxb0ZyQyatAb3OQc2Wyrebi4a67X8DhjRFELoh4lKMRunOHUqB1VDr0hhYAICQ/ier5Qg7BhtIU
6N1J3cSZiPs0/pV8uNGi16sjQSbBU6QNKMKGgXcMvdrDbMPkC6x8TpnJFFmcGj19++jdnxe2Uyom
gyS8mlk35xQ2HKRm+Uw4aP9ncb3eLdMz8OD3chJxOMVwYEoq/JvKzxfS1zX1Xw8Y3nNcy8NGyX4v
pg4jlzxbiGDNdOCbsQRXgGfoRCaMAiJi3xjWBad8z0ageL2dZkmDdHFqd2WfP6jZ2pgclFw0iDyY
t8a54ffslhcFlP06omJ94e9gilfDGfhcJmamuWmBgdBoVTMQJMDqyutcCISADKvq5IVsOXrmIHWc
elqeb4H9g0Fl0WP5ousoKeN0TFFU/RASJTPbX2tzifQX9VEs+b4NAUaCH2UvEM9XY0JSRWtInuj9
Ev9Rv4p+/OdWOlEoWR0IqDg+1dAXsZWq7idqwL3yp0dm6LroPp0trF1UEdIbq/kF/rjBFtaM5z8x
70ILNpjNSLisVvcyVTbQOIyFtHvwZrB6DNiuZplueyy+VLEUKmtGQkFIeyZI3SRGvofCu3OJf79N
R4BOwNlw/vePkfXrzDPmho/3zC5lB0tMcFYtSuA4TMmxmeeP8a0IZ+MZjoY6UeueUENee4B+kmAM
5oL56xLRLH/rttTlD1RodYGSupxHiu6prCS6+lkFfV/6nJhi0PYAbvwDBjTC2Fas2NJuBvi+5bZr
3bV3trg1FR7EykChmPiKKJXwfgJX6KjjZ/KIWTeG/hzt6md948IlAwbilE7s5q1EAtfpEG1zapCY
U2eaCSeMqYC1E/lzj0L1u1+Oh5dlCG70blCD3a8/ocaZno4RZBHVn4xg2znwYx5UbKbo/YzJcLBu
Tj3ncTnqVvkFme6hQOudA6T6RTliSuF7r4afcXrfMXkgCFp6DERniajeqNe5fmn4tC5s1J25Laoc
8LBUnec+93UGovxVSRxXZj5wj36Wq1r7DZV76BQKQXebKioMTayEhLHO1qEJnM7DGhuEuzn9ZhD7
FT86JBRO/zJZiE/iL4LrlG99x2/59klGjwks1gZf4u3X3a8OXSIQ7VRTASx4yXwREg8iiPMhxZFp
Hl3UAHRzxr9R37FD68ZOOxukyXaSMsvarFJujSTqr60uamJRNcDnAW/uv8zPfmSfpbNjxHHZiiAl
ABFy2b24nYtdQRPw89U5XYjZAIjNb0opK3wVpqITHA4716DWG+dWxAEmpp5dsv02PH+Bu21+W3sL
08mtQgfCjJHbQJtdZ0dz1wORX+NnDKklJGtql7OdyODSrtWjU32xO9NMyvtRsH6PnxpvhHdR0qI6
YZIl+ngdQiS+sR9DJyp6SGjW0s7TBPfLO7u7OBv53di9Nn8HbPIo1kgRN6/Pv2MSSdWIFlno5UPF
8F2tiUm0Z3vDBTkaF536GBubydf27Wgo4lTC0dsXsP+RRtXpWR4NJTHz+DgtNfyPw3TPvnNmsqKL
h/v7pCq7utERLq12CMQSE86f3crvhTzdIgFgMs6vFeYpD2ZcIQxQ4A1Nqhsv85DIE3/kLKM+Bbca
GWYRoUW5CfsAe0me4qQlkekNC/kle2HEagdsqHlU++cFR9HP/gEVBJgLi6emyWIf2isMk++7MHFy
6ywN50ow1PtTbWovamQVtF75VUUckIPTgRFDpkYQttYvtfTAKqE66BpA5a3FkyRuPcraY9Uk1R/i
R80hvA2orCXJP+7HRaURvBvHORSje2a7VWRJHtXVSwXJ/KynIUfQfugzVxpuKmo11PLOpdx6kCZs
wDVChoR0CvHr/i+yXO2VvGqZfJaYQHHCdKH/eEUmYmopbSfU88b2jsbBoe03VdPx9dFaMD1RANir
KROBkD+AD00WfcOVNbbsUgMONSd8BixiaMOFUAy/G2dr3NtFuRjk89zYFJhkfPEiNmAq/INXZ5Io
+cW5Nhm7f1rkSmEw2o3im0uYMpElZhFijDO0zEtFU/4dAA/Tgm6gNu9/2zsueXD2s9ajRWF4/g6j
o6Z1Wj4gemnkCcsSQU/fJKgZpMKl/Jg2z3QUOkgFyBQYoQpMvHVQwh0Yd2ehHQcxlLskLS0H2o6E
bDvtNT7M9V0MyP6sQtrnK5tgZnCh1q5+4w2JRh/deO/tN/J2by/QbtKPLVTy9GA6bNQC+nD9P271
Oqjci353ekmXjrMDqqqKi5fkEE3UDuUfh+bmyvBKlO/2xvoTrnkUQSFvKLx7qX4KE6A+uimcPqgf
AYEvy7A6w4WdTxvXRbOVwqUmGeJN6I/n3DpZd2tfGQsKbGu7iEeacqlBAs4ZECmzr8R/iAW3h5NV
83zNvBGGGvdrJv3A0hGUO1Bk8h/xwKXA4CqJzwzWSOwo7rD76qyG8T7kbA6V2KCThrBMk5YE/g0v
1ek2zwb2KWqdCaHc0INNAY5amPNyiIa8G/7ggGivyDZRQU6UJJ0ygLgVh/t8+byGiWJcJ76q1fCD
zUMxtO348B1+E2M9M3vMN4GQpIZ82VrO0TZuPxwzaAQTER+PuKZEAsEBpUUg+7nnj6uIZhQ28/kG
1cjBVlefF7jh57Yj5xYz8p9x0xYfzMvB9MXH2L8HYU7Ug+iiH/Cuog4RkZK4wdDVts+8XKPPfbxW
iilWOxZIum17H0yB8PdgAHCLrdPMnoBDZVWhhwFCNlMV04vOog7RVPK5W/PYg+/daqmSDXYOPH73
OPreDWiwqumjvSUC8PUJeAimvbRy5d74ylACjUc4bABaQY6SrHLzC9XmiGhyqtYnSC8YN0Q1t8BK
lAIywnXsUNQsVt+Ep5mQKWt0irpnAm22Vn6PuexFlqxK0d3HmnVeaEYLq6rZXIaPCKbMYlttAfSr
zUJ7pB6FXwVgRfNUzL9Rel/xzR2CUZXHWlYkjPvJXC/U6WFjHX2ThsYjVGVW324VGw66l7e86mFa
w9LhyoB0GZgjo3hFzl+ZXeFfmWEAgvZBJ0wkyeLkBY1wPoX4MYYuMxPGEsbcN+SS78UsEtcQ86x+
cEEjEgkjD0osnA+JiAIUUa4HLpdoVZZJL3TMuGJfSKpPJk+OPpUVQx2e8iokjjQbzIuazTogD5ZH
Lc9QU+Xj9nNuFxhcWPWJSh9Ku21f7Dr/lA1q6+zPvlLxHJUKQA+3Xk+n4wqX+GyGHLLXF6AA9Df9
DGUz9GYfMytDbsPprcJbW68EMlA+g2Du8lagD7/UaNih735o3tUgHW0x95gB+EdEFhHs40i+ytGB
mP/8/+Dik+t2dq456kCVTvDmyKBvgRkVgmzOsPvxY4ehvnzuhVBnmOvYktHPFR4F+v9PZQvXuFDc
H5vM1qfZhnREZuPreIbu5PLAhOFnzi67f2U4UojUgQSaKBQkOk28TCuyMOjuQffmy2TAHrVisvXH
g6X8sHLI1rvC5Yja0Ydtsos99NBRnHy9/EKJJkiaEYVmgVkOMUrlKPd+IDDSu62j7lqbGqyTTilg
rHSOhQJ3c0Vq/Gtt/dk0SNVm7Zp3DjrerjSAyR3zH7CsWvTqgLSmWLf9k1LgsSWlaDDx7duHUShK
42itLgRcIZYlpMggHKsYLX3qAWwWkBIrV+n+MJL+6ghPA3hNBVZ+ygNfmZU+Cg9K7WNfS/MqOcUF
SQ6Kbx8jFnGX1JyCuV9xRs/UiVisvCqHQMc5t2puAUN63epRjvrdnLtwhrk87InQ08q+84/rovlU
5UpeVO6axcW6oMOvMQQkvrIcM98hSeOnCM0U3ah4FyKVqx4hT7JLsAAR6j1uNQAqtFeX2C8E1rs1
tTnbTla+TzUWA8SJ180hD3rch5JIZ5fakIsxvQEzGVNWOucv+jcBY66HvyudSYBuhNsirB0I1bnO
y3vFRyUpSzmhO4wwd7XiKqq3I4EjtQUQ5Jk6TQDzUH9Eqq5JMRuw54JWzytPcq9Kt97A3vxTS1CK
d0NOitx/oAUGJN4Khd6CvYUkLhKNEZpXf7OtHQsyV3TDq7/nQV/rovVj3wx8Uzmsuyak/t1gl8t6
XhzvIt5nEQjsvRuFTTHjQd4tOHqG33G+CfLKE0rcpVji7M+8pad5DNJfR/v48uxpzLbt5hxKund5
HnLAImPehgLKmoYVvDUn83coz80IZZ6Tkq43fMGLJaVFhyhDxreNq5j/xeaIfgM0odreZTUBsm1V
fyBo2r+N3uosT00jIuQjf9FYtLBShxVuZdqpY21KlM2yxHrlOYb6yAAcNxK9dLv8+yBkQLQd+3Mw
xPClS9to55aoZFPz/JLzF99eUgy9pWaRfDIJb2FAOxhN7C+M6Md0ziQALA03oKShzwIbbuP7Ff/y
q+AGZDOu/2XQBgMupeZMYnDjpqLXKzncvuCr8iatCaZ2Kl+xvM1KPwh/fwWxVHR3IRU0ukJfC6nv
THSOvvrc6bi1WJpmWutRa4ohHMIxx5YXoVWssWnfP65/A2VKAFijWeCnK9hnSr1ic6Gu3U0oDm80
B/+62AurRTicHU/tfMvx2VUZITGmK22yAlmWJrN+R4DmFm9CC8AGDqfnSSpY8TTx2JUvZ+u5gyNl
vQzz0IWzDj2gYllIh9T3UEKcv6vUb9zNHKL5bV8q29S6GugUtpwWkOHA8v1ALcMbtfGOkYE3e3+I
1dTYqLIYMxXRoE57jlyHej24GkrxwrumzP/c0jSGQL2rVfKqGGDIHcns306K0/zxFvJUYM/2cOon
qpx2uclGfeii3mXcgCnym7jui5WxOBKuF60Ko3D70EwXhRMEm7MhCKORgXlVXvQi0EzLvvL79ZIV
TyBmql5d17KJJUYR2aq9/ThER2SQsyOuPwcQI+1nypGEhThhduZeKoeG/cAJ/1uYLt00ZYLXoPTn
i2oiopQ7HAZYoLnNHB6yaqjLzX4JLlZWjUxsSamNfohL1zB3O7S32ukKE9y0NM1MCmvRrARsSygZ
qUTgrArvfkLoguguRJ8PJAdRHQmtAsXZ2BGQ8X6l4ogP8Wo5pTt0mDNYb48T7o1ELFd2UfaREQwQ
FADP65Coy8vz1xDCXqIbzgdisPitQ0BAj6mD/kzv2roq/yVWvC4Bunt1XyE609oEwof3XoZBR268
r+EdVp9BJI7vIncVUtZK6u7TKExqTnj1nsg/nKmAuft7GvTZ9d/L4eznB9NPcQ95AvNmFodZBJGG
5gfvi8zOlOtMJYXhjA0a5Wqd0mwKHclCdyzoArQYlUHdARc9UkwI8MbOwzYsrip11GTe2euFSovu
HjHW/P0K2omFscj2ezWtdK2qk1l1EdL7VqWB05a9ULW6sKTUkw/FjSQBA8GfYEjfNQBrCCuHehYa
lDv8pSuFCS04jrEDVpeeGDQex7Ud2/AtfxcPT3v9Uy7Rnm2VJlvQqNH9VTgiM1SmzvRDDoye/eCN
R7/kFS3pMMA2Dui+x4PaUGwSJf9GGkpJP0OsxFpRDvepg5mlvnJDFgH/PehkJcT33iQ6AVz9nCpT
6JRf9p6CQylq050riaEu2b7KB78w3OajfJLlkLRYfMtQvvlcLnja4gQ1aImp4BM0iFN6Rge/4uzT
oH5lc2MO+SWtvoMIu45WirXEMEB+Y3aSx3mALbvTWgl6cWzCdJt1k4hbxY+uQE+MTUdJ8snrb2m+
Fj8GJm9rfs29YiFJZGTqbt4MMoFWbyeGDGGdyy4TpiNTajcj2Bs8HQlPJ74g1Nls78QcR2hHIQgo
R/8eaI40uJU2RV1oydyACs/lA9BtpIkdN8HOx08LBXIRGm9qu0Sso46LkC8p1hR5vdp2SSX2XRAm
XmQvfbe4xEwBMNK1zwjWaeYWF15JoUy0c9ZkUPzqDlHYAd5U2cIoLkxrvI6G/jnO1lf++qTG4VO5
XKCBnz8+I+AvkSPWSOLYyxr2x+iB2QB8odJyIyejCjMYcD7PBjcroKqLvFejJWBwnnuqYRTbGWYO
hAE7Lq7P2lzzNGz7cJ9xxrgMsx8f/27k871imMLPrpNJATDTXHpXj8QYDiotA9qMs3SBWiurycY6
GARQ7Ar21hHEWuWAL7mCdXtyeaiXYm+bLRa0mOOsZ3rWYKILmOga5soaaYdmpuGvnFn7ZjKxVqSn
nzQixicgWDxQbWJ9DDbssBIiq5b7c8jtEidoQ4IB2F1xpy24ij2OhJGOgQKwam4+wgdRTHNDNaSO
P27WR95ypvNmwRAK9pRyWiXV4+2VgZffYYGT016cRAJhagFYGP8VjR0k/68vDT8tEVb3K+qnO+uw
/ZCkJGUF1UTD994M8T+XfzvmpL9sXFuENG7rGSUiqXlxpt6M54Tqpt3cEbxWpV4f6dF7hyna53tg
dO26mEdsjwyRi/aAwPAsmEbRsofZrCFksCDgUA4f17AtFTZkf7butlF8YCCFzOV4JNglKIA0ptCp
FszHT2sLxish2tYGVqKnf9iINAlCB/AfCkCslB1ARhs2gyux13Sovwp39663huOw9mn3We5t1Aiw
NgcWC9UGOFcK2pcQfHwE/Le1vsp3wN+b9SGE7IK9DBB8jvtsbziHVNbQW8K9fzvP/MM61S78k+MR
Tvm+7TDBMX1LuG0oq0yXXAuTsgIqcYMVvN8TBS2Ds5pfa+79koFEW5evN7yX2Isu+K06utDQzoQq
758Kd7kJ1to0vHeNEnk6Usi8TGJ8IFKLH9aiC1C3icU7zHxURIs60CHVi2zbb9QZreRbBWHa6V37
TTEGmZMNkgz4OdvLU5GCBD6kF841TQx0S7ok+15XzyB79Fv80FKtQouH/ZkcxndmniWqbNxOyupi
EMoj96xMVv3CtMmLn0e5vxpkg2NEs52jYLDZJAFQWSI72d/VE8ptzt1Ex394z4Puv/T5zhlM1O+g
FYTmjZCjdDGC/CUCyjka2cvcuTYIleD4HTcrVT0ZGgTZlWUwD87ii4QVSJYPrBfmWkjbMS7kgwdn
tIekqir1br2BdO1+GWa9f7WR7twSSH4QyK4oOcESbnZq+qwsTPiiAq7/bU5cb0KiHFsKlZZNNnTt
8fX1nViLYbFPptj5qgoDx0soZ7wZnD37ZTjdX+Jma08aV4JerMULsvC/FrNJLP2l+wc1cCzv7IVj
Y2PgdsKztwXAWBfkUPgq4gggth665F3/iPxBTt0N7fAyQ6Oz0wHjgv2kqt0dOPpwhQfQFFG8t9O+
Hopn8rIgV4zIOAwhl2xJ+BFk81nxEgiE07JaAKWSuO6nqqYsTLdQOv73eiNeju3bNBuQRsbK3q9Y
7/zWjOUuJDEXw2wMm9NJXx1jqPhN8Q6RdctTrN7AnnZJYD/Jr9i25WfMMdmXScI4sRokE9goDpvO
7PfWJt4dCthBDSAGVUeXwygFBxqcYgrKY2ZRjxTy68OtpCLAuNqKuDsJVffbEqhJlQAH4G0H/H1e
Vw9sBbtcCM7t0nztYEuEL+5zFTao88uBt8snm8Jd6YPNscqdd+d1qnValng1n+nAQxMAwCYr9WTs
Okk0HU81MigGl7oqPfiDWSttJ+rWccfY3NcUbhP+VBRh73huIeml93v/pl9xoF29f7mlNvT3/LVm
zoquWj+nHnbC8hWBL+ACVUN/SrTK6KwF09m6Yp6YLqUXMEHpAoJUlurlWC9tB3oUdUONsNrm7sjx
8pHqBdKJkBwGFnfzPWyZgvMpVJzczyTqjFm8s1wqmv5jZtC6ZNkXOSNjGkHAH8oH7ywZFY6RCQm3
CsoFljYyhsLooJtZBiEAMmHcHCkU/mP4bCw0amHWri/sMzGKSa/W8LJ/8umjHjYu//SxReHRTGxt
0ewmoapxSPnBJvxhTKG4eAFhkqumA2r9QQ5MyJNPoYLmdm3sbJpNcm1S84VNaMW7ptfUkVme5kkI
BzJLbW1H4CHuG7tI4etTruV0gima+rh/p0yL1lWxLk7/9FXfubtP27z2tIwVsnGvIPZ6iemMYcDL
wa7P7a8Ya8Dnvk2En0EgDZWQWhiAB/FPc59rldiV2lV6zrH++cYt6JOGgGu+9CKKUFO2T1fwPPEg
1dRibRy7rANw1PisPqyZ5HN5RNCFeXnQ/b81wSiqvUw21qVuOGrmw9x78B6q93JO2A+j7+zsV9U8
itbBV9AxVlBeuGXogp/bMI24ubhutlu63hBk9seHudSQb3pY1mlGN4QRKkF288QB1jCBtQRkEcuX
HNkaYgRT0jPwcLVXwIamtSCHlHP74pt6iSXv7SfqNkOiZt8hR8IOClfTnusevUXMhAb6ynP1kuOe
EZWOGywLm+pusERohSHDUr/N9lOFgZBHInE9WqXxGndAMsjvq7Sphq9EiUC4yf0aVj+rXVDDJI5I
Q2O/RBo0NEME0yOi3W7Y3EqAMygeO1wFgU28FOJdveVRzNTkM7Yg6B5bomPxoYHizi2R82w2p7hd
4rD4F3Oy5PFk3KGv4y6gS6MDV+H4fLD3gb44Y4J4XFtOTv2GcWRehymArlrveGj6fayPQra3D8j8
6MnRlwkXx7MpDKmQ9m+5YFdAGzt22RpdVnKNwNWyecJRP8s9I0u6hgsv4Jk+0JWc/JpeGizfXAub
MfWJFUTOAcabLvqMxIxrtCbhMJnGcgnlT50FoOyp4EoN2mmtYz/3aizY/ad+Hy2M+IxVyHI8YfOB
cImKjQld9Td4NRoyHuJTM12BltVz/Lz6GNEUvDKaM+fRDvofTGROktmeAjJAau55p0IRguqUY1dt
Rng0T42r244o1cMuM/b4cfS6wQYeHi3gkRLuH6FIoSo4P/U+o/4d/Xsy9T453+fSCQ1t/Jr0AL/A
2Yk+/otnjPxRC0zS0I4gyVOFh6O06CWexZdUml70MXZDYvPLamu/SWSFN+EB6S2IM+wTdQqMBfoE
e4Uyc9cylaDAmHjaAbwVo6cyb17TpgKBmplEzYQ57gk8ZGHxYxRSphAqc9CU4/qWByOjhytlXFLz
N6EjixVXfk4DwsXgCkHcpI9g1aTZesXBidqzWE7oCASIFrcVaeiWlbyeGJ40NsunFwJbw9Q5+JP2
GMvC1xBUWPxxU4rUdQxuLVy1Vp1r5f2zIM2JpbWMW/eaXJcrQjQlUdimcjcr7/8q6Rw+xGVkYsqv
JFdU5sXNCMoxguED21IlDWK8Sa6v/dI6x57kXTIWtmLAwaMtL+1Q/ntcRU0A+Ihc8hFPnMgnqYEG
TghRoXWWi2ir735zfRue2QrznajFKu2jo0kiULx2WXB+xz54I4x00FYqMj+wVwUPDc6cxUwhddZu
hlM6A30p2EDouzwdtcqGwwZsexQ40NEnDNoPvn9Td2+q0NH0NWUlSYbOG6/suOI+vtDx4hZF6ypA
CEJ1izBsVjSYgIeelBhdebMc56Ks0U7wzhv312Paj9IfqrW1Ee/WqGKMUvk2r1hCkvMiq/KJnkbm
DO491riBPyHP6SWIE/tYjcoRC8gbvnij2sYHEcDUm8V0bx4QVb2kqaEPb4k0ZbLBvFQ3k2kz4oF2
PSWrVB0xYsdkapYe+TOQNlltElTLI194CYIRJMRqDOAOcCsTzQfLmd4hgI+73ngt0SE4uW7IGETR
5foDu0zBsf+2lsergRLBMnKG1BKzapqj+d4tLQnUm3HoPnwsBGng9U6C6zIS6k/gnO1yChZAux4e
vDb1evecIows2nSgRLxKG5bidPzh3OymqeQIXWv/F5oBwk2CQGqbUeqcubzn4++Fpuv0CkELLns3
Aqubwpp7jz6nPaQJFNLQt5urvUoejtbSQNvPwrUT7HLkMGjcbp8ebmlxXYeW7zT0FE+XRjCfItYJ
lnwEMlLSTVt2nmI06EVIzw1jIMpIM6tFi2Ez8KUlchBn7aRiCfvoZKc/hvwEhJ/Oc2Nf6Kp+9TPU
GR+ZvYPkwP0lx6D99Ccf9yppZ6kehpaA0e+j3iMxZET79QcQs32a0yMGB1va8ghoYzww8vTCJi3I
cJmlM+tSMQlz7mBj+0kTdL4mNRIa4QlRarYIFiRMQTJ3DK9IRyU8vj/yNOwQRpge5YML1/oEtmkI
LVzPycGIhf/Y3DPpffw6lT2TIao9rNiriyGv/6HScVaXDGxRpvy4aN8uJpm0DKwPGBjtYEW8LDGZ
t91OQ9hy/DjFfIBKeR7zL4sp0iZmDvDezBSihz/hlDV1CiwOKkVvpoC2W7GxzPkdXcAY1feNOaO5
TazAA1nixHLHt8rx0gR3VG/EtWYhQy3Oen52LG2VYTn+nG3BKv+xTlIVDpBJ8nRf+EPLtLX6tWq8
Z+JktWHSJOkdRzLZerQOq8VOEZ43GfITcAd89ZFTJYOuh9zjksG0sjSspvq7rs6PNVIniX8OK00+
L3WF2mZiyME3KuHPhXSt1wPIYxN4UgFzR0TS0tcs2YNZgeTiwovYZ8FFniKgT1FMeSGNmDEwtU2h
3l6W1TaB2mqTBHh2GzX+levOJtUXRUx/kJsc3meillxgBbL3Sbcxv5UD8D5vF1j4xG58ZaxE6j3l
rrrmM305EW7d5KOw5fx4qF25+QK26VQxWQmpeh2Sx8OZZPwa0f9kBxBKaveKkdX/MvdhbhrPns2J
AjBmN6hKQw17/1dbmyZIHnaqLNFWO+vtEnKM0WbjOSTZxX6009T5g7KLIXF6SoxZqbzV1ceyycDg
WpqR47anZ/xUOBDogy4Bi3WokNXXmM4hIb34UEDxd0lJHS9u9FFmlsNwh9/7JwnnCvWG4ClVjsTz
iKWMYJTJm+CoHmDt5jV7RxLljkI1Q5oyKMhGGxgf3wE8RnOdQN2VEE758sqrD339o3G0LUR+7r8K
b4KaEMcQJQrco8u6ECzpcrg1tyDmPzRBsQ54T2+CppTTQSycgF4AGxG7wVpAfTMVmc7FT0+lFo9o
aFsVD73+Yp8SFfMimds1FzyGuLwfRSG2EPUi3J7Ns/NUPESNMD210egIe9TA+wMzv3nMj1Vmdz+T
hCDx2LIXWOhymnodpmn2Jd0ZfqaXw4OP/Rl9xL6ixmnOaqx9NYd2lZ/+7VjOO7FcK52O/yxY25bv
RO0NjQuhZOddD5yG6q7Fm3Hrc9KmvDQzxMBpxcP73WO5gdeLRzVJwt2WLQetneDlUV3ITYaXIv18
2u1kTIh/2fhD69TCJIpN7I1q1jdqHPw6F9sC6iv0sxNKKPhnkvd/40Cp+trWHI5e4tQc9m5JB8Az
rOCwwGKEdwMMsynUS2uUr5qEZs2Lsza2mbGD9V3UlVZmWypNm9g825PW1af29ZVibuI02SYCz3Bn
/XFNZtlw5EHXa0W3X2tPMejkEF2jyeVFP0k31kzjV/kNGh34eAqbVDzVHs4lPp+zOO76M9keerAl
vp8OXwNNbwvNyQBRTjKSYdMFNIhrHEn3xpX0RDY6NxK4tHWPKSSqr7dRwcnWXWdDXiofmwCAy/a/
n8L2BhVTwJcvibxwPl6EZao4NOQgsgPmVTL0U9DE5Eti9WHkMBkXeC/XpswK0akTdpttb6QUy472
04qzHVZX/tvDOpPvYvzWC8DzH+V5dsxqsWQLPgry+77BsQW4S5eolWa4P902/E5KchlqL4ljBmzW
YPDy1eXXsAGDJxPWQArfGkOKH+s99CaoxTGgAbo5ozlj1IyAkamCquJxq5E+q6M6EYL/vH2Su7h7
FXrDKk/af/wq8Jxjmi9+15gp6lPulz564msvuv5IFpVuUulbFKaC/K6281930efysKlf0z5QLAWP
PsUf+fH6eNkFVlPmK2tFPQGUALM2XE0d4vYsFBnfLBXWofcedO/AKsfZ827sDRjdYnCnXXQCpGO1
3TYysQ7r37l0jJs+SP62URX1QTApPpdM2Qr48g6LjqWaMa/zv/q6vmRhqfOYixUq6kHvdYjMeXPX
WzeVlYPe7FVSe/D9S/pti3fvQQTIUHSAhFHqYZA03Zstlzj1SJjSTpgMlSQtzVBf7iI+yHlnH8p+
+G7WWrLwr4WPotLIREQ6SEhD4FfPwQfZerEl5xVK/zyKkzCdREsFEZP9ezh4LE6Sl7J1aSviY1Qd
FOKFg1E2woCX0dab6gLM2ee9dIj7RSuv5bx07FRJ/7kD1tJPZqyjcm7whdmY4e+hYhjcb2SXgN/E
54u1SitOuo1q57ouFxbfcfZ9PSGlAtc5E/N22keeIib+kyF94BU6a2LxLk2U1hxHkvsc9teyC2F/
d6MYHVWQgp9sPKw07ZqwDh1XlA9Qzckk1HootdemqS6VkbavQEeXaEDRSYUKTFkYY3KVv0aVtDG8
c5k1abOulzB5r5wbqGSwo9XNSdjwmtTSGvkKi0PAj40gg3E7wuZTyNqL8KarrVGvAP4hP0XM+Z3C
jZ0A1MOnpLA/YducWoPkCkHr5dLDeZxcWk6QgXhxdDk34d0ZiPMYCZyunOshBFuloyNfeXTKfbxR
mHpSjk9nuhwHj7o2ezonC258KP3kOAEAM+WWXzSmbKV6E1Qvn3Ru1IcqMWh0jEXO8Qy84IPiJi+O
psyRFpX/bhxi1B6HozqyaOSdP6mKQbplEf0mEFu7qboFsq8oIBsCJ7GLc8lRaDIiGjEb2Zy5mQcw
56tNN8VjsokWv29g9t8Nb5CRnVd7M0NqKw4rZ1XIjCkIGrCeyUbtqeiCGce1g4gkf7XNQVJ4CQGa
MIb9LfguZtjcffR6F6UJ0mm057ZH/dwNGzsKePE6rXiJ9X4mj5wvMLGOZsr3aO6HN/8/J3gBuwSZ
/6np6g+g8Cd5AyWunpShCMhpePbn8t3KAa/ouOqeyGR+vhKoayFyrb7ieeqJgiMPtIP/zeH/F7p/
nTYV9FgM9CCxigP2sBs+wFiE51Rmq4LcdrSZm4lT4Gv5QGySxuEIr+LYN0XoGbr6aWt0WcCpRPGw
+gtNyL5oNcRs10cFksUbubRPqitcXWJr2fljKQbKFmPoCBCYqcpBr0p6o8DYLJYqqMHTvUsdSyI8
xjVAc/8pmBwIWe8Y//pu8Gt3DyIXspCQd/0uE2qyo5AwGV7N9oOi6sD8+pv52K9m2dZjaNGi+xMr
iG79BHycde7JB/oU7hNfvNfL+vW9XIJ4Z81vAIeBiTpxaOS16AyhY0tR5wbMs8ejqHuouftB98yw
rtQjkIi68rKtDcPthXlAH52BE4gKisX17tpMEOFudkeGfkAvNXZunh2MhjsGCa/t/VqsKBGZvHLW
KqQ4dLFTHJ7WUQ8Qz/o9r6DF1xhX77ZWX+U3ZZKO6SJw9bwZcGTu7nBX9NukZfw2zC/yqzs6U3GM
RBnaAFMpefJH5W9sWOssxgO5T1sR64IoALcxY79GGZX0tRvWSXpFPcONqwGj6NFHQ4S+TCzAHJVz
8Inr+eRByzji6BYD3w71/zwrdznBxhqLwC7g5PFciHsAxlrNeQqCXXjrJ6ugIZu4LYhhs5h48wj1
PJcUr9C8jNsV/KbpwXe+dGMAnMzQM7U+9yWgruYixRQI2ru9+0NpLX8WR1hY0fA40jqxAReScwhL
OnpVvEEfBbTp0168N7276rrKRcxo20Cy7GfoQ4Gah4awTBsrjwp1+OTgXn1OsqIVDYXLHn3neOFB
K5VQShpF0tkrix9J/E036hLlhLt1VeC/220H44peNAG7aFGDmEWx3LSdChHWZ3OjJfKQqD9jz7aL
r2I4r67j/omA0pIxLhVYkJQo6daC340mhAtyWZrqL4S6KqBqVNX/LpQ+HBGDJsvohppplV1bcxH/
/9oSH191DHnQNx/KmwJGRNdz+7Rv4G472pOpnj8OPH3JtUTN7r2HMdj0Aiw5d+yIDVuhRhettVR+
tLvkL1UZPctomMP4QJjg0S9FBO01KlgN3H7HoapgZGxIMILAkPkZxzh3c8+IQ8kAf6hxegPOQVI0
x8tZJ0xENnf8oM57MO7z0SokXPsDJjz16SZuC7HqsxteZLVawyybeQx70Y+Iyeoc3jXI8TilQTGl
Y67j0+MVRsTkEPy9Hgt3jEfnlZcB2jXmtLK0WcS4mNwpgyAkXmaC0q/fA/jhf/bXaMHEmM36lFsT
v+AqiVPOnlvdpaj/4PC9qPXyPPVkRvF9IreWAhwxWjc2tKFZqQx/BS+XEdwOWhQG+AghaLT8Okrz
3Jz+X/fGMOjtBWXaVnvX1lGlfayPfjuQqlCEUDvgjbbX+qx5hL8aO5L6r0kKrkMJWJoEIdce9RGU
aUbEOyehhPWOCCPoypSE+OuqaEuhADw6uWuLokwsUCDxSFiq+swU50imftJbNYbM/2vkZ8kjZ9Tx
G18wns3RyWoR6Hfugitw9kG9vDGAIYsP/wHOvx7LTdseQ3NcaUdGLqNZPsty3NqfI4mBNp96Alwk
DR0pk74VWBo43OEzpVW/UV8CE60ocS00pL03s5IPIM/Z+kR2haa8x9oA4fsaX7+YDlPWgtCPlefd
LvT5bR9V+ZImh+qTaYlBakymf+i0AyzofeCmrPo7KZtfeN8SWI1j3Qi5DtHhTYLlKHVxR8DY+YJB
BbR2BWgPWAhUFt5Zo5WSeoKQ0veEyqgRiHEczLLJoO1GDg4ysBu2moWIZrT7i9vfQSwCkGw0B6bf
K/lQ7JVSjGi8bAzkW3fNDwOTCrbvkdZX5k+nOuIsDOI94lCTwDsb290xFyOc2PMdi/zPtrDTC7gL
w7SCl84mZktrrXWWzXEXz+tf1nR1seaRqCjhcvyVfKOyBB7cJb+IproyktUQpCabm/kS0z1QRXec
zsVkkjAJKNytVlqFZnoFvPTQdiiULalVGz3V1iawjxGUcUjY+YSlbjPHAp/aCrJhzxhgJ6b7gml6
RNY5eYF0xufqolT+XPSKeMQ1NN59yEsh+LMEyjMA0bT8OMLcrYNwqat177jLUXEpYTkgHfC6EQVS
wIRS9acc7r9XxXoIcfq8sZ9q3eYnCdtjGfcWe2k1+k7q2KPpQdCThQj6U2esx2qkgDlshKWYtTIM
osgYvN28bNt4GBn7nJk7bA5K4cDAE884k2se4ApbmFjRZEW92sOMWhMtKNWDhCOksjsk5gBswreb
0NeCgz6JggFJ8i27Op00hYJQcOLUwOS2A6QIA2kUel6f/eXNm6ItJMAVFLyK6GoVgrruazlW0vFG
/CY6K3P/n4tsY6NYt3fqaviIQg+rlhZvb9R4Vtmbjyn3j2cXOCbG6mvSeWbSXnn72oUgpsUZkInr
rW69Mw970JiE7QqmuY+GOKgjsDc8byx9SEFWbJk3JKnKi7/Wz+8oCfq2W8e1EkU89dEB9jTGdyDX
cbxo5HkcqN9awfj8A68yHZt9yQzZj/j+aVKmXzvR8YJwI2kPokynlqsOLA0zQbVjgM1nsVa+8uQY
7KNSr4H6EfEu5wEacv7Tdt3998f7euBWgjEWdFk8t7jNni6Hp4dlk1FE/VD8faK77MpUdUMcSFqH
8wLwOyGYMPC8+CILXuxaVxM6lCGDIm38W1G+o67J99t++wrV2SILMbIPFalxePUOI0nbezJmkROZ
augJYnQ/pBOsNtQol1LOoQ0lXTahmwRefuUmHNaWwACtdvLxhuwKQCxHMOF2kKtlIzXIxO13cCxD
0CGotYxPExYK7QwAPupBV47YVt9gmLDSfHbiztITslFESIsXRhBC3a4PNCgRbKSpXR8OUPZtJ82x
VZ9usWsROKiKbHJijyHZXyxS+ZtVaunDLN5j9sXBQulPC4v/hOZI9x0zU5mB0r04CjMOosqpSurv
zhVNXZkhBOc+2PnyaApRQRRM3TrARrpoN/5nELw+poeIOX8hnr5kG0dHlPxfZH9qPUPWPF6dec4+
tqP0HPXQuEhUREXWUozveAo0fLU/np3QvWogHM00cYAdbphVIc3Yt1BaA+cgZ6CnZyxnsvGShcz6
5cL1DehwsIN1laYIaf7MLttVjU+uaYHawxlQNXK/fHJAtfQJYJ+dCekSASxgK+wV3iOVaCz1fe6t
DwGTGJoRq0QchKMzvkDRFTk0x04PE9CCxPn0QOT0Ue2KOjMC24uIK519gNS7gYsl0H8oe9/9afh/
mUEA6Ccr/8tj/1t2Rg+C2D0dFqZ5hnG/HaTryP6cBVYfT+fbg+oGGBG2JqIiA/TibxA/WR8N81yy
gpqXBon3VSFk1mK0dbI+LI2YmWNBxr9dUdVM/tZDFucKbn+ETqZurr2NKhoOKnAG1n3PIZtXPggn
tx6vVvV1xwPQ+VKvwON0rPq4vMRPD5XiXGDNsw6vN2/DOveVtOTD8RcAY1B3hv0cJcnQXWk8JG6H
7sjexaDx6xIKgHo1lUkX22ub7QfAJf1hrCszvci5CUOkaNRPPksgso4NzKWW46f+ZTzJzr6/goHa
IwOdPGcxaO686Zk6kr0rMYPInvXD34BOhZF79yeCVBBa42qjZqxx+CaLjqzllHWdrCBn/iFVertw
ZS6sLjLCHOebpW1Th/tQJMrByCNafv49z0gRbSM2k0CDNfGkSi73ST6esr+n2Cy2SLswt5tHAnqJ
2Q5oNJNT+d8rVjVRQ1D6abH/1Z0FEMRrIWjJ+k1JipbC0/jRj+4lOPz/w2HNMoeT7pZq1FGBbas5
oLzrT4qNUpYkVGEEgUaVhRrWnUz3vHkYY92HDX0VsQWGdrj4PAhBa3Q6QUOrX3xBDjwID0c1f4RS
VDfZGLyD94AAI6mTVg8EEeEOSs+ZNXld55aDAZzV98s2RMhrRrGgxMegdjX6+9Agy9QFmrTlI4lI
1cGibbu/ByIuv+c0txrift0EosrrKocxkJbnBecX5QvzV3X1GiWUFivjhnIeiFqDCCar12EeHNc+
YGmwR2fC6y3ij7mjyDf+7mV3demXkSmqJyqF8M8clTDevg7a8F5g8rpp3v1xmgnOnTzGFgvDDC1Y
EWL3V6Xm30BUyki48RqKIONewAFOdvLtdk7ibneL7P4qIkCLCJwmPHNiNAddmTSzJPjrlROxvckQ
ucxPh/BAiVId8r2330pf7Z32FtiIvVW96gZJMatFKi8A83B+NS4B32gAD38RVio+7Q+0PIYTZf4X
EfwCdnOHaweWrxf3FeLv9fBR+gQNz165J08hnnIPmqyDaeZB/EvUPD3VNuBLD1nW0cEpN0KsNCVg
wY3zkcyrmacPrOiuVxhAch5JzIyxDuE9db/GpoPn6eCKfPLwi9RvdwUyL6PvysZdlAtTTHryGdEv
H9qDpXVSVrbJDSF2sPHsBDmwgnTDFOCTRDhuce0k1vKRmEdyAURx4kazgcqdSgsonGuf80FevyTI
XCNRR0WglFCPVkEXf0g38aotuRdYZk19bxx/FPpE/TFIz7QvpgrSVcZg195RMpAAEELckJ7o03v+
RrKY1NMXZtGs+w/dk2Vulp+tO24tA8MJeb69ze72upUB34f4hhrlk45STXaMkBjIEWN3Vbe2NEP6
ANVCdG3cN4qEmNgIV21joUY5BUunDPVH7DMkuU2XYfkSa80yvFsk99vglbHmC5v5wPEBOQYymx+s
BvCDCqS3TXe0Ku/MAYzxM9Zd7JekQQy6rD3uQa+m0F9SVlrM0SOxvcsDP+PwvsS1CxoVPoGWGh37
fKL7xg7+4gZ+yhtxZu5ygZCM3VnmdH48BEyk1BurNWsk5HswPFpUQ6HaGkuWPJwguiOMApQdNbTH
bpuBYxaPjQUBKftQ1xYkrsqL5Uz1KYvRC1xmEzg4l0sxhsdSA14MxgwAj4QmzvFDBwVhcWn+IyDB
Kc+nRCBufgz2/YG+A3mqbvncDqOfSdq9+gUDZRkbsF3VFCx/wljiZSoCS66McnG+4Ys0CTTMNRyf
1sI9l/oqkmD8y5e4TbxPwf/r0Kb0ZR3NeP+wUl3dngJOp7D9OWpX2HAggBaA8tNnZGLXCCXsfP/V
SUmXaId3hOIrm6efnDzjOUxczRLxA+saIkVMI3LC4VqE9GBNHk8taLD326Nqlh/4uSpJMJKAzKpE
5ft2dB9LlJy9J03ggj++Ew9ntN2V8nSM2/irRhYGKRycONXZ8JYPqKSNOcfovmyDN+07Ou8FRMky
CexbduSRZ4vZTgCXxsrPbxIKtCKJQO2H3z9o2W7Evynjph4XzxSNUlgvGmA8TMWWruMwzJpk96x8
cZcZf/JCHeXmkdwNz+wTpg39YREZUuC6RdzSOzsM7LeA6VsgL8wESSHjfcrFSq73HOMkxmOVlm5h
WkveuEvIcEgvSc0XMecJXllwjXjz/XSQsAjOG4fuXi3J/dY6BOg4ZyUL25BYAU7O0f3iFv3w2ILE
fA5V3bZWtAkQAEUps3SDKiXA1vB1428P2cjO5mpmaqtZ41JVDXC5ILHBvwaG+ZwUrNIovMIxaia4
WWvQ4g8XImUVvXlF7IN2UYRCi2bCX9ZqJxDjnr6ahAjXY/Ib0CI81aqWto0r51odjkQcHd5zDe95
Uuzog7GTGR3inJSsqFO3ykG7+ZHlazTjUZbmzPh4b/I19YpDkwPkPYFGmHyhYMkHdBPvPlI/nwgP
IpDYaZV2YYJGvbp0njpEk56RxdGQH1wQksXkSvPj/QWP2zndT+oDndh6cF/6LW9tvbzuXp3fV13u
VAl4ZH9KrH4uDjrM5X2OtvyD1wI5kZsP/ikU6ZivQhq3mEIhJhse+i0pFvn9S+KRz1Z8uU5F/duN
SUhT2YEBHRDPiCkvpNVPQt6ZjWeBRuGQWM9jQNjjlypjWmb5OibuPssc/N1NNZqoOE56rkDv3JMR
uge9LEd/C7L5idfHvSd2/9BLU6g7eaTKw2BKpmx5CX1CdWSy3kqfYl+t+u4DtcHKxn07hSPf39YJ
7nfZOkqHrFuzzY5jGms1C59Xp96HXXu+E12OAKApHEs434KLuNKbadO4QdNNbQCj43yVE/VJIGbZ
KwTNSXgLFyLoRBioAmi0+VqOBzDQSaN6s8bKPGBAzdzDB8bU8WpyKEJTgLocqYcqcSp0GWZMbWBp
WKbnPvhBJd9NjdzjJ8Sf4LtTTMckJGUiufsioxmKA76tB9lCSHKDMz6o5WJZ5sonlgG7ydswzHeP
ONO/hUicQX8xldSFXEmn52k7iR8G9P73GnJAHn3KcOoLAMwoCQ9ejzwRQCbITE8ev6lwEzteWQY1
lQV2Lf0dmO3e+NROjQj66/HwW1W/eYDmGpqb4SBhuYpkM96g6Iy7dCDvLDOq4bl9o9n+mVIz/jD1
7jBHwnZ+hGWhOA8p8xOp2vatln6vntz3fqwUNB/r+Qwg4rqhf6Eg0ZlFjmj12XAUZcJavydcoTCQ
LGKjbAIKMgDyr75TsqfB1bz8vUw/MKhu0Unyw+DMVUHGfq7XGJUpbjWSmFc0R7EYFfVxPG9ldWLe
38A3J88MEnFUxBnc3/cV+dQyd+R2fJNULflmJsKwage3296mVkvsZKgL8OgrYj7wLODRTODFaKRI
KtJhhFHnUnY9PyQTt6uBWbC2HepmX19bD70kZcjDuPGqxd7H8JKl11Lj+nFbZnJR8mGrG87KFUpp
QHLaazmTJXgyQH25LbzqINzBk7dF7gByWF52rcb81wg876sYExQWSn/ts1tQTSn4i7DBUyGNJePS
vQ0cPZQZZnQ56G9fg3wc052UfiLBvjdQcTnVLzxa6POysyA/mWDIvpYA9De+QwElNQu+yYMA7mAs
ve1u7HR/hlmXX49XsFV8FMrpSmE3gIktF4Vq70pDGcdIocHgErRqRqDERxViZshHstzsxthX+UvL
tXP/H3NoXTnhr+2oL11Zx9jZ9RgA1pLYbmFVJYfWQjs58++QKxdekCNBVpa9jZol6EZnJPUv1xnU
yQmEQQh7ASgGau7Jv4tsTXxrEu3GsnjAW/STzKbQVBudi2j04TgrHejsL6ngpTaqzVs+VxXC8uqh
WetxkQbImIhIUtnF9bC8z7Qy9vJC7umTfbL2GdeVNfZmJmGWZDTAMpVxTfw/jgyN0kuDzJDsteNk
Qj/W2Xq6eL7/ePDOMMXjzlOlokOb+Xt1nCxpnS9/ZLMFOj3NY96Ifgm1BbMob3DcDl2xgigtIDxF
TdhhU0mBFT3HwsTmZEnsz9xvI41f6/a0sps1ceQWbdBLDLJs4viljoS8EvM0mgjBNyh5BlxRwRzk
M7zAUqIbEy7tApZvg5+/XHRYZ0jLl2o8cKL/rMbqfPCDuTZgC/5clhcDLKfEG6kPBipmz325wDWd
xGBP0tNojr7zWZheBdvqoeiXFVgSEcExhcZEYX/E+qV84mgkOV/kv1+/aKNW4oCBlUteYkwjwFKG
WwuBiNuXtN+h4eAUs9HT5T2pLUwVBKAwVNDJ7ICWXUqDnQzJRi8rdraUa8acf74RnM2junBLs52C
aMksS89l3iPz7B4rutnG1Ph3X6GB3MlNTuhFtARfI8FinCvLvwWU2gGMz9diGKU5vtAbUUA7h3Ij
HAs6j0xf+smB5Hex9e3sRMuJD9z7QqPf7kfBzk8MLHu8OhtioSLiXSr3vfGkrGDAX36f53kPRG8H
HKL2vf4ms+oVvUDn30SeeP5wQJsD6kvN4EWUOFYJV0cCAA7iyxEuzivCzaIPOfl+aWC7yWaERvUT
4Sygu/mOGQIPuIntIwrAwYRrQnGdC5ZM+iMKhrVlWPUkn9ohWmtP9c8qhcXy8ITIaa8MFQGtoYI7
C78KqHYFlWuFOaLRDWYNxDz7vRSKyg+QYlW29Ow1lv5Xr6jwg2+ucSZZdnqQhbrLOl0LsVzkaOMJ
T1YrDCp60oAaIBpqwHsin1FsGQUjxPA8Ywf4Q9NaoscX6FG2wzqoMUxML+MMIAEODttMr/KVx2YV
DaBIz52B/ictIvWa/dzzsp/yZx1x2Pe+jasWOb3wc2dW0OM3XVbPapZLIc6STdsbToR4vHEmtu5i
I1wH5Ng6ReUkWAsCDxn63jWJg+gcuB+kR5zFs/rMu3mExrmSvtfCNwicYIM2PAU43XNGq9a+kHgb
T1Z7LXxrxgYTHoZJvlsj8IIqKyvVqs9RJ4ldDw6RTpfDywTDYPLsShgFldhKJXYdrE0u4qM/oFbs
Tv10SrHdxtRO4sMaw3rgdxseTohqalUAYpK5V7OUWqWpPePrrX/2hZ4tw9SFITEBdchrd5FZxccE
zEh3me/17Q8NayK1da8GXdlWRhVCdPgcbeRd+rL8qy5VC8srn7VYivBf8Iwm3CTxYwtuI4/7mwJe
lHrqxQJw2uT/jVxmisUZswy9YyB5kapvKqpZvVHe2bc2Wrft+t4Wu5kIfiIuBKeUzwfKq72bOSD9
Kb2Bgs5gu6P/5pJdqHoC7M7MxO3TNNCCZQrtbZVMrb7lgSJS0ljdFnjvD46lMR5BApDkREHBrP7n
ZyvaWxTpRm7OzgyJZZmjruwf8wr58EjdecyRQ0Vwf1yf94z9Pga7cTFPqKrK9iH1uWoz9W0SL1S1
+UOHKpiDMZ8GD5DpD9dzMaJ6LwWpHymEPy/bKFt1sINiwIfiUca/IiPgxnXqB7wAmLFnstVIEMhZ
cuxx43kzbhHUVpmnAT1wbzLBN8vmlTHpbZQ4M960B/Up53+LC4nkAO0uwC3YPvJFrYx6D1frbo4C
5u99uetema5kDMLb1MzRgSj5zVGEVb2XX/O/QE+YM/K9OoZUMzknv7DWm/dGeaqbNnkeCBSlCM7f
fWVEFR7UHu++JzBRCqXoUBY2QQOa4b2DuZxk8jdYZW0QbPpWXrPfqVZwlfDTm1nme7xPs3pMEAY0
4b9nF5mhv5D1lYOUY1ktIBR2xAUJFK7uhwvRTdH63Y2iZ3DcICN75irT4EqlS2kmVVygjdqLddKX
sbDDmA7y7QxQpJ1wJmgs5A2zdHO2GOKaTi+EpRh8qSxugaTpP+c0vddzmVimxx8+djUTOb3Qqqdr
iLdTlM2h9WSg3Dp436gc2U0M1ZOmcJJdXJmGEcRyiqqM+YU4/UjnSzrbd4Cm/Nv2AyzzWjndB1GH
nu7ky+AKkoMQeSJy2Gxr2lGJVR1JbTiHGgAKOMIZPgbDdRmLZa37GBwqeDetdbJ+Ki1fwHtsF9s4
Bg0tc8cCaf57gJEW5BEtrUTFqJGUvwNMeSQBwZXR8yrGCG+3F6J9XFKhMiJG2HC434GmF/86mA84
O02d9pN+psH2FaIZgkVJeUEIz4dlGZiRlBLxfQ8D6HUJIUmp/SRmdRfxiO4KXqY0tmtvuqWfU/Rw
ho46QxNxVKYerYIaCoCGU+KHlQ9B70ro9JkQEI23uGZsG4rKuPAS/vxJmEJFU6JGJ78Ss02c4bhD
IdugKHn3PhyRoezLuRKJ6LMzNu07DNlDT7lXJUQNizK0cAyokS9xSjniCQM9X2aiUd48UF5Q1iHb
kur0g/3th3U5v6pyLDVqUaAjNs+c5La3iB7ILhvjVBMFhS0CvxWjDlEIycmo8I5ebeVh75FUxUCU
tmPQ/jaZd8GJ6rb2UeEufwJ2KXqgdi4ceDJV26j22pnWZXn9y0mkiezA2U5bOxtS8WEuYGRbjsC4
czi1c4e4nWFybAXCk9gX8lFZnY6OFgGVOtYdhXj/JLOsKQDg2OuIcicwcQzyQr5Npq6jsaSUxnXW
aWzk3cVnpLbQDres/7GHjNHF3pTN2LmFy+zKVKoAs1hXs+HZyoNFBAmFhkADrSx+znRG8hGp2wIf
SoVHCggf5L8Vc0iNm5oTVjPSGcoO+1tuGdSm1JcuLXdeL1jfseccdnKqkWLV2X20XH1H+uXvkauN
YUUSOvlN2bye7gVTMsbKhjlsxd5C4m8NCyofpY2QkHAFunaZUYi9XWxcil/XLd3AIVfwQyVrWYKW
EF7N6ZxgQpx2qydyqciWUUMJBvRuOKv7vKooaw/bjFs2unEwwJbJLS06v4qVeVwZQw45zYn8Pd21
8dJ81ARPlKegupLMFgSdnAMD8NsjL4WQzw9mpjH7tEBv1RYnZicw8zfULVYHuDaGi3+NXPIdgupE
H9pPzKy/hGUbepUDbYht1ott+VLyJ6LAHEE6d4LwKjh75srBDmau6yjS3/N+U1kmlO8Pqj7D/mpK
PGL5REwC/mu6uwNWSH1g4R+XtKU20gM4kkumUomRJFi9k6XOLcm18QT6knfeP0ewVheoa2/SdtK+
2nJBpw5UpJeSYALwe9Xdf3Jwn3cnh0hWJA1sQvziHWN7ImxUv4uNGQHrHZokdNrYaoabaaMGc83o
5VdLdS5tgZUclLUEyC+XPQSZw+fSDYdss7urLlfN40rbcrj6/HWYqZBdLQuVJ7SH/aHPMwVRgBuL
yPGRETpXcga091qJyDcq/0NZ+SK6vNl/uXBfvRA17XdCQX5UVY+izEBheIqcItNApeLetuEs+lvE
TRoVy4xBMsFTI1wqOeLmWkmEKFpQFKRZ5yN/jXeIkvg5vFBiVfraPO/DokY2iCAhJR4P9LGnqUzl
1FZhotYyd59qSDxxUVU6TbPElppZcK/RuZ+ZA8iq1j8SvrLAyrVk1B1LAT2zt6NQgQMdNoFDATwu
cGTlxLtQOHmcSa4AaEauu83UjK7WT79mub3U05v0ZQBbQTamFnUL2snV4uoUTolA/2aSamZVBAo6
lWikioMH4mOzfTrc6CH96dadT0SbSZvOHuPRQ0n4o5CvW56Aalm9NSRa4j8d1ENhnTT8R+Fuheml
9kqNjW3WlLsh8M+9oH3WPzFG2aZoXUciKiQOSRCmsmyBjxs4B74T28LZjg7t4JXHUfgvpw7hRDUv
VzIiFoJLKtz4mvg6+NVcNsHIN+6i0FPpANPxah8zEcaWI8FMT+fqGdFukIPT4EklJOtAHKRnNJGV
wykhnVPZvcRJJ1TK/b96ZXd411OQr60eCXKEHrp1yT4Wu/mkUpaPj3+eU0S4l8l0aVKqNPuZloys
VjrgoUZ9T3Tv9tUzBspT2G07klKrv4bTKFKqXRdI9YGP/4555ByJ1ikcAhUT/E/Bk94jxLfGlu2w
rf7IjqCWRaKC+SbSISYheEaGiCE0y2frmnM7eZc8EVPGG+VMsi5PTX1YVupiwtzANlifiHUkVAuz
SotdweQXNth2xwB9/A4g/eg1QlLaV54CVvju01lMexjB1N/DQwNfwYEWcdJTsD81OExShECZ+0PT
8xe9ohZd+yI2kpLlwPQUKpLZkSj76+83VEyqt/oYZT6ilkGGiFwWYB39zd2/CexZduQg+toBpH0u
fW8r3jCmL4nnm6qFKsIm44nszhRa4FgTBrTJjphQXX/Zfw0p0KsegVzcYchgWiO3tGxQ3ZueZNFg
q4VF9DxlNNgqDTBrycz4V/OVSyf/DZmR2T9Jc2L3b23dxSowHYZcN97serqw941ZBBv+oiXMkWxW
edtG7ifVHgJqzSq4bYyxhAEcaeg38jXT6Wf5GgHzSzjalIE6Sa6A75CHtAVMCMXZyP7qlKIlC7sg
OVq/HUg3/krhCPtn6MX19YlUC6vYS5yFe9UmhH0vc4VcVdW/4/Xz/bu23yv5i+KF+JiREpfFjQKW
gIMs3u2BJlSud1jV7S13bdfjghOZEi19U3MZdNeMPzemcpfOmYpyt0Whkbp0dcDMsHdZUCNl64w6
I+/NDoro3z/r4P6XM4rvaR//8tfpORfBkBcwbBVjiYXMlloG/Q4o12XGH4Xy/lbIrAsrYc1qu/0W
K1iegwyhAvA038AgV5YlaJpIF1kyFElQDHUqVgp4edK+FTrMO5hMWdAzy4681UWV+0KV78YstFG1
tfRBOZXyLBXU+my2ylmnvSydM144CYovbwGhWlV7AhJo6sGXXivzov4TysknbXjRGiEsllukCK1L
AxBg82F1LHGgqDjackfLCy+Z1bOVMrvzu3s8QVmmn2x38LfNhrZS6O57eAEqlnnbtph0KoPy93Sx
pUQqE7QFmk88ai6wDkMypB3V/a2Hw94DvO7UGYlMR4EW+zBpOoM88p/SheD53aviMIanCIeqVl1G
6MuMkakNMopD7zjU4bRnus2MWCrlcn7FPMMjrq/d/eMBbTkDa38ivW9LuJH7d56z1Kd+b2VcSssu
XcpFU5U6jE1V79jhTHZLKz8nhTz4HXRDfKyW1yBMBLGqrSpSill41c4SzoOJ52sZ+qvIDHt7n7dy
G/T0QyZpfXO5f3CdBJjDEnknBmnfDCCxiRvY+BKh8tXYY+4osk+6diPNqueozhJGi5wb4gAX2KHM
YkuJsK1b7l0wEnB7CrRcjnQsxRYaWafgiN8YDC2ffKtDihu1kGNEABNMgyRJtwaw5Q8lZQU6AP4L
PZGw5IL/iW1mKNI13s3omVk40uc414QA9vjTgZBxyibMy5IBO6A/lDxwh9oLUnX46hVl/9suwFqA
CVnrZysN8x2WFowiVcU8+UUXihJOzAQa3DntHa+KV+YA8TAzpmn0ndHnIFddPenRYlUSA6HhUhCK
YYBPIg4gF1Bd9u+RpN2Xwbr/l1gkI1OKEalgwbRCf5eGUoHT5DshcaHF+JHksAiozWgaD5EIE91b
VLTBXabjDEfKV6c3Ho9Hu0CPCIatzHx83qKUtc3p2Q1VF0nFrF+NXc2iUkjiOWfhe3f2dTRxEN6j
JPHMT7MMcLjg6z2OEkbDnzwxEMUZtgXYG4iS43Gz5MmjLpaW5EjFefXhAgHvlB2i9guivL7KxM/A
diF9XHvEiJlsIsO2VVugzXlcKTsTN/aFzmU353ttsRr3gb7bRJxU55Vzo+jOAkj/5WtoxZkid7BT
bFODs/dj8g2P0rxE5KRjEUFXL552FcuGRTdhILZLpBgMYVD+ptyGv0g7JeOoBBgsyZ+EME4CK5B6
P8NKOBnEkdgcaGNsAiUlaHyQD//vHugIIq/1BK7Bw/1JNlNYHVU940gB3OFom80ops2/hEchmp0P
3AG0jT9HB8DCaHr+pxEfwnZLuNwvrsqMJ9dItRHU18r7YZZcN63ydknLRLZ0MA2SEcarT7MyMcH1
+i/nbV4VLfQ0Cwk3UGGf1aKX9VanQOjwystcZywKLtHhvd2DkKrW75uwvStif+7EIxUrmlvOeKEG
A/XSRvWCTAs/pcbrFRQv+j7FxOTPHLkNPPILqBj7S2zl1BudFdP3o7Z8UpbxTsOE5jqFa8QceZsF
jCNr4PBf/vxbu8uJBEXdXq/2kYSWCPmnq1dOs1NeQ4w7/TdCTqnC/ybrZ7YIntnz5tgUNxWnGybQ
RMt9bbyIDhjBDQjpccvOwka334yLd8blq4jZqWU2uMnKtujPL/DjKIUFaNrsDaJs3xRY1fCvr29W
zINcvv4AAS1xETdpyrOmXo5+jmmKzTju27tkHb5jP7ydVo9A7YgR1/6tQ9nd9dTrN6yWTCyZhUnl
qoGn4jx88WfEGu4XYgqSobKYv4kvjxkLID6t5SH3GMoM+Pqc2x4kcfMzGIL191y+LjjLEnGzbpKF
UVGbiWf4baqqjh/tdqJEcYxESk1zsj23fSYAZ3IhkNwgVzdVGB1FRDF07/xf1tmCs8z/Egj74Tyw
Wl5T2ABNvJG9gyHCEPgeyCEVbV2GLE50PzOPQv9AjvKgogSBD0/KqaazChVAbCmg7Fh+l6SoG8b2
uVhfBpAXVDeDLkC8Qc2lOhLNw14esgeIP24Z9nH5abgIH5SFd6S+TRl/AMDOJYr2ulTY+GLRS041
mOZtk7NUHX6VVm1QPqhnFNwAjIG3lTHJ2I7gXXYme4piVoBP2KuSsDSXdIckRdqIueoVViUK+FRk
3ioPLQZrcnexmMiVIUj+XeNyZvMiHdQLiNH596IMrPaC+t10xXHU5QzIqnR4ABBUH2xsy3m8FWLI
yO9XlLCoihWLbMGlU/EeHldjNUUsOowYYljHqHaQz+8e0igKH1QH326VjeYPjye1FZVTBF+Oq8vj
EBtW0NLRMhCrHstw0F6r5Rfu9EmmgISdzKLmcr6TBgNq+TBGQ+YLxt2AcqdvSYqxrYLo2EUbRESd
NmzPDLOfa3K/uhPC/e6uzs/H0X6K5mmTpLGPkYMVijPSk6R/wF/BcsRYne6uCc9JFSb1OiCWz8ie
KjwSSzeXmTZjGeBJoNnWHuFlMX1U7zvxWzem1UGTh0Mugk/JU3LSCXR5bRHrb4ohqY257wEwLdrh
K/iUtSWllZ1ipIG4SF3fZdMHyT8AfIl4lTgVV9yxaWxGxKw9cDxl8OkzihpgG+ylsktzn8Z+77xD
4Mac+23ZFd22m+uRaBPur7CB6OjQ+dp0AWUrUvv/PHwqzx31ZLzCNqeMRzMuww6Nh3zVOJ7X9/SM
2nqE+ldjg94Gh3ywKRMJ+iuJ2SRKfDmiTzQwOGsxZWizeYIGawlhNRClip4A9EGrCcPe84GGCQVF
7WizUf7Y/ZqkqGZIWngbz6ba4zlSWrKUwfwE4AFU7npEaBkOuCDctM0/ycqZb3ZfQ8B/smY+qt8l
8RKVX5tW4+Q1SzzOKgUs4lnE4XBF4c20JmXEH/Tu8ETDTaL1dD8iwzaNxC36jec0a8cwWksckRpR
jB9apgMm2aTDR4cvLHxmtJOxLabHiICy8+nKFgqo2+u63ciPpRzIw7K3avebRQ1kLOZE82KJdwR+
5ZKkU06As5YtCWPmTeUIM7Z9K2+ILTuEmtpFDvUR1PA/m4PEr5N7kTbYtqGmrztmcjZSKhaDMPHl
/fvuGcX0BO/bbMqZPXkL4OLzI6pt/oodtdgt1amBYtYqHaDm0ZxmNLdFdx2L659AhyVRCU+cfPeY
yo1fczC1OyUHi4H80O2DUiVomY4pFSyuje27Ln73I6TImBxIGydfMilmXi7vJpdkQQnhvj6e4OxB
ndmS818noUO+G14mTeDbmUAMeBlrQB3iPgAeOwpGTWQma1JJG2i4M+rr6tMhqPNoogQaIZq5vz2u
eF20vOclhmiRA5kARmcEpxJq0vRYakP1TRYZY7A/1mnZhoZGv7P1DJ4WjIzLcYmgH/ayYuSFHqXv
bPpSSpFwcIlLzNmdRzPs7a/k3/sJMGmjBUgw+Yb0B+rVt7vEy4DZFDuhewSXHRPw2xIhw04gpkZZ
XVJQKgWyvAD+DFkkkaligqq5GH7yFoiBHm0jOgJ8/46hZavyDfkASlUPiRTWQ4zUK9zlHX/2cOwC
pKZPaQAG3doen58Wf8ZZJkh2pq1JIuYzmfZroQ8v37d9Lf+mGI7xWqPmwYBGlDK0P2LC4P/4TOti
TPAJdpSwL7m0RZPnBxKuoUUJAHASjJavVdXi3/gxo4lUZ6rIJb9KD8wSjDqC6M/CLhw54NVlZJ3E
A46r62+8gQ65vte/x4JSnJkMBFD4wrtvytiFUpygU2OERRG+cBQ070UHPTsEHMnz64Hn9FAVdWO4
5+c3U8MAgNwln7KSogLEMfJLsrPG3EAK6YQXpA8X0vBgIu+myOVNpRyJIsBfnu9tdqs52lnEuQxZ
ufyRkYRLB1cAymsUrlJrBnmCwfXoveozJuN7v0ebGWFSNmv9xxuMlEcoy5OpBHR8l5h3FoIQUIwX
ZPfHpsNyFXjQ9PWxI7WWCjrRz4rF/kQkALW7SkekVyQp2Rwlfob+IHjMQ/AgzSQovFqdtr/iVW2X
nvA+uMQ7EamiJxh/1hXAW4+SLdzAXM/BwCAxq8xE7cpMoUpIzOVFp0lVfDXiD0ENkIA9/5AkBl4a
SHFXuxj+w3XdXG31noiGiImR7jd9H7Ff2Ld92g1Yc184aQ4ngkDtbNnpJN/pBEa7GpYtSv+aztsO
tXlWbnZefnkYp23nMH41LOsweZqmu/3UyUxIlq5xDIHwPvATLYJbWqvhjv2mKLZ6AydHkuAx/sB9
6ctNgdZ0SIr0jqzPPefpaV0QP+iwgb9usGyKyGIAa5gnnPeXLL8lv29jk5QrKDceuaGqVF7HZrLG
WETln8EFQyva9p7LnzfmB8CUjSafXi6lAySDk3DWate8XuM/HRKuK8Ow7kPt4wPpxguDMGrR2FPx
bznQ703w+zCGHJB1fOTJV3s/n+fw0z0WpWgXR72ivAuyXFGetTP1XPJGCuKSgyuvV/xkrkHfxzs4
E0I2Pu9JvrIRTuBJkTq0wylzsKOEfE1FOGnW/FTiK4gdvbBBSqlItqkO7hHLlkOFAoVxW5/Pldwf
knSKPoL8eVLrqOYSmcMAjow4P9JYN0GtN77CDA0naGFeqXHf1jAQO4er2+LLjwSRfvbqH76LKO4c
LAQH+84VcxO2av7eynMP++7J8Q8d7Nl8UiwV40tRUVxQpj/+oQpH8QrzO1M+jGRDLMj7QbCBDTqG
/tNjCM/ZrSFc6ALED543NeMt6yAsVrsmoyoKyMoClTPZFUswT/zvtcbouDvOHUhHlblEgdDV2t31
AM1sjziB2GQdWdWWx8F4aF91FFtCvN1a5foyrvw/Im4/zjlGSnJwvqP9k8AKZ6sp+jMFWlqGXk3T
QG1iGDDvJVOTj80RI809rF2+lXFy8JPkVOZf/fooCGa6f6S9enPwZm064ePCebwgdcc1A1HZ9VYm
S0eZjf1vU7tzxBPxS9Tk+8p6+nkMwbudZ9j96y1maq0QdeIg9duw/zdD+HyV5jB4q8Z1OuNCk6p3
GyXRNsoMev4T5se+C+t/jiCgRbZaEQLnZK3mPyIzlykUGCbdSkANC0pwd8U+ELVpWFNBTp+ByQk2
8TmPXGtNyGalSsGfjh6eZCMlLx8t6Ty+Aoal28K6sI0OEtw+uysGwxFUBv0/YcglT2KCjPePXSht
4MkuBMQie9hK4n9H+tmxyL1bkcIwj1C2iIPOWnrlWwhXwLJ9zclFI/yhqVXoDssRp0Zdm52cXP88
vxjb42yPIEfBeRvSSpLp8qXCpYg1xyFqRh1DPOq1vk4KG2W2LXs5fd0ldw/6GHWcf1Q/12wAFrCn
YZDMYL5x0THPxAUqANxjXx6/rj48gry9YIDmKQDTVZVrim2YS9z6suWsuXn9V6P2teeTyg6Tuofe
M3BR5mWLe4yc0VHjCGPdD1Psol2lKmcilhcf+HCDVkLmTTcS6nzjVnQbslt10hnvfnd6A3l9unAf
wdZh+mpVXW0BTRVct2Bz/UHlwjnMNFZSXArzMDhg/4yoQD3750CApoWA3zu89rb9ttwPplwFgJm9
RK+cTq1doauVwme2ZT8dzWQL7gBtZxxdV8jt05dHnkWs/x+VqpM25VwF9UZ6kI/FqBUsm3CiKN4X
GzF9bQPDo2Bx/vgBUbgEl7TZ7/k40gIQVu4KZ1xxfFZd0Fa3q6V4pS6LpKH//zT9ZnvYRzr26iXo
np33OiMLaMBnKdgCG6N2yke/9auXCeIXXm+jU+wxA+kHl2c9ePcsZ6AeI9AfNqtzPES90ZKskxNp
7zxfsP4j7Gq9epgP+/1IMW5FEjqrvmTeE0lVw5ItHVfmfH17U9EYCzghMlSyT5AtAb382OpZ8lRk
puqMBgL32Ytd6zODQ5aIBvWXBw+Qaz4zjOSji2res83iNR6CJmztKKoUAExULL21x1GKf03dbWxW
cTRmy84oNx8anD//eZly70isawxpA0uKwWifwdxiUwQ/f7ren9+0/xXyoaNDN+B3wfnE68ccu+qf
YTkt/XBd7CMDQRNl9lYPHiZDqXYS/s6JqRqMzDeQ9JxqAzVCfkEqKRlh1CJor2JeU5cTKbq+8txV
ESPwGao2qXY9V4rj86KzLbg2cSYZ/NDORFISEwSkpdaCnJDUvmwifOE5FLB490lJypHR8HYD8grJ
jWlX8eKmZ6qj2GVy81JSM08b2tJO02rEiDwkMS1v1X2URSNUPCo8b89TbIoh0uHkrugpO63S6ZoI
BTdjAwsDoHrjZQc5F0ehLeoMa0mGJhs0dvXHos3Vo4O+3rTTxw6TBLmGh3vTrYr40gNw7qNoNx/F
VMtWsfDGEC9lBseJ4BCf5glwamO75lThY4wm6HvFK+Bl3hODW4mOJ8C3NkrRc4IFzUS51vpqhJSi
nsoQwnt7oLWqSIoQGnRUbvNsbqqvVHtiycqv4WQTdp2CmTLRUERu0cKpp71WWHgmCBA4QSO7YUAV
G+quNiP6gNLvK3UwwrSHubBHk2pMkdBxVIOQJvuNDi4AMWzxJbSCctYuS2fwGzMzZAxyJf0vW09A
0L2evaqKqyo4C6mzcNPJJnX+jgo9a1zOfoCEgFetKOG8bKL7KtAdDDlf7mQo/L1IRhjIh4cPLNdP
Gb+U/B4yOFEAZKypbZIYF+fp+gHw+i2Uvhre1kFWV90blDP4XUngISEmJA4VUzqXaqNvTSVfEnod
g46TDl8NbYvx+CFvbill1lVUr1IlwsP/2fVOrE5OxZBZwCpGC+GCUAiKOzwPcbCP35JmHh+4PNSN
D2o4BJh7/kbrvbvwbgHnH3xZfVimMt/w9of+imgDh/DE/rf2oq6JM+KSN/OAeH5f/HT72q6wQ/dL
f7Vs2dR69MjSEB0FF3D/QEfxl4wL6QYa41s7Sp3IGw+BaeIHj6rddsBGeo456aIl/y8+A435RnxZ
a7cJjFAWLZbTJhFDn1ADDnzrRCLMXiLwU8PglZ4h1B+JKGA6M3dSrhzMIrInpPWf/AxvTc/Iafvy
3/wxF+5sRPAL9dQuepti7HoA4vrUjW79XsPt1xEvEkIGl4YXBy68E64l3QOWpa+ZO6AM5dSZ5mxp
q+nmKZwNJihoLrGVzDVaz2yvFgngGQsC3XoKc88uD08tCmkfVuVvjColgrvm5pUfBvajXbk+bvFO
mNKA6PhUxrNn/xYhNLeD5eK3BxFIWg4oQttt0Rp43u4DQcwMqIdtzw5KiZFyqZ2EsZXAclfXAQER
L6oQWBdAIXCN3HXw8bViwCFN1T/QnS805pFYCm+zzX6MxcoxGah60e2y9xn50wmxzCwbaXwm1uSN
YLO1WCDj7INPnSffTfk0vxSE4mJvKPk1LHSOKX5AGQmphCFPqyjDlG9vCWFUcFARQ0F1jZMJ6wCH
MF9UJKLFirVRNwt8mb0yuB8BR7axDlhfRB7xJpr23TJkIPbOFRZ69Wzsin1hd39Ingpvz1Sy1vO+
/v2jv/iQpJArrpWe8E+a2ctyL6MzvVA0qq8YqR5WhmW4U/XPYnSORO5RwaTGYktGMx+LcjfmbBi4
EdCsAvJBKlSmGwOtDsZNXDn1pKnton5S+GBONYfqNHLgoIeFkQINVnkVmRXY0lILeM6T1zTxJLRL
MBdSo3EAcPT6CRPRnJW5l6bjGj9/3ljX5ilbjp/A30Hklasa5pLzyg8egncKLNhkUdCIWjahDQdj
Z3LYbv3SEkJ8BUdyLoDQl9tYce8wtJyASWCO8NvwBEYR2Sc/y7KrEPQqE5crTtaBWLJ/0lJuUvcE
OchNFGov8e8AAowTHquFHhP8XV/b44TcRF9/pCcvJ95CPCWZlTwJm5NbFTCgWYYJN+8d/YNE457o
5qBOXPsOsUPDSAB3/rSE1WQV279HGMnm+63EJcyxkY1ZvBmnzYZui1ifbjs/seGFQDGZXHSXUqK4
g5Aiwq7Y9QOwI7fwa81WY+FPjLY5OmWlpe40Iggh5e2ZH/PI0NxYXDeL+8myDNsLF42fdwZ2LSW+
joIqIZDQ7AiQamtdFPMhEIzxKc+QBb+pMeWpgKtZGiuLQxytX7ZwxjPnfPE4YSZDYbnF01Dagvul
1kOsscEBnhJLgjEnsMC26a7MoToUT9XRbamv21BFJP1YfLlYMJ/rgKrSniGuZ8yLQdscW7oPx6ex
xlkTemHEwh8eaQXq3eS9O2kyVODVQofvSkW6IEUkSQo7M8XWxh8EKW2hJE8c8+oL2cyFeHklPEWc
7y2t19Q2wlBDpvxSktg1BPZuAhvFENgMnnXNVgeeZnRcWHUV+Yk29quXf19RHtvqZumL4CzDhzkg
vzM3mJajDaAFZqCYGb5ktQ/yJ/VEqNOkGW8NMdUl7SrN7joZjDnNvDEvO5fMib2yY2lfiFIc9a7o
tWKs1Ht1lSW7+K8PtZ/tK3Ww5rg5z74ElK3g5L/r+LN4Bx+kolOe0rUpCjwh7SsKJQENsKDSw3X2
b28ybVzmuG9VYvRgS3ygfmwWYdYlC0KBi7+/ISCVXIc1c+XL63w8gxFZZGMjdQnZk2l8uDChw7Dc
Pg5vL1GSwYkL+T4TT/gGjlI2BgPiAcflQebooKAZE2R6LIP+w+DlUHFURYebIAQMzxGmo4LvBE0J
VG3xEHUzhq1WhjahIRnTdsmjmPbrd1qNSPqVs9wV2+KjR/1or4Le9XlgPygZpJa7l3U8YVFKjPeF
IpGNbwYB0+OanVjpFT+5uxU1joxti1bOpj9WFQXiIQ2PkLj4mk1lrwKEzy94cliB6m2Qt78JTkpb
U3YH/sk9oM0Th06FeN9hsbhZuL8Bl5rceOzZbbU+OKqzVtnJu7GNRZckM+5Gg/Pjf3JjqEn3909j
f5xzkjgCqPomyHbAmS+gIZzpbzrkrvC9383USBCOXd2zme28olSMI+P/VGy0rS9fnvZG9F2C6md6
T0opozd7xpybNLoi/YlE8BRLW+5vW7p2gkTttdmjmBCRL7FLWoP++gwPLQkZQ4V0Z4VSxFPdxdZW
XwdPsloP/xiSsp7W0Rb2i0l+DAuuFd2uB8j+GSykf1/Ra3s5lcF3kdXgFaoVAsyHjKiYk7YdUGCX
PvazWeCUPqZFD7+efNfLsokiN+az4sDFpIeTCRSWjeHMYCXLqw7Sg5DD/a8RlUO3yVH8OIqUfJ11
rOMHoLBrKQvKOyywtTb2HuxmQdZR2up6VPe56tMSntSf1pKCnkvouaSagfgAS/vxY5FX/oR8/w4e
YMDm95XQ0rp4krgoMF6PIYhJEKsGRPRQ5Y3xR+nV2I1v6n7IZBDj10KcCaHH/lACKfM5Myjr0CTG
2XN9qceJb7gD4Feqb0fJNXcxDuudpFWx70sb+NrpIlJuhMQ8EDsQt6k3fNlcryNDfkkstveWn/Id
OCtI7JcEWCnKM8hreqlrNh3zl+yiaTF/c8xTBP5Hxm5VenEbtHpmqPBUOHUfooXu23jlG8MnyZ/b
L6dDQfm0FgqzTdAEe8z4AXB9iCQQ/eMYymDwot/McEC68unA2HsCvgfWAMZiPo+zz3Yfx5mz0c2K
GVrSRJ+1ns0a2lrdwlGpKn721hfGnk0+Z5BlOG48HD5fNlLc3cwMUWov1dmlDhPDkbXnaM1hrrc8
Z1//1qnA1Jj08MytqFRb7c/Gzto22O4V3kEG2KlvaoyFo22IV8hbWEIlgJV8aFcLgm010G9ANlEX
D8ynriGD7UiraGY0Ss+qCj/A03BlQV5yRdnXxQBKLCoZgSPN6M6BL/m6yCMZpGLcJ8O8knwQhw0r
E1fgaSyuRHPwbx34iYw1iavhcl82suRfbGIFF5VClbmSblsqBp8+8se1ulnEepzWZrM1Xgc04WKj
/PFQYu6Rtdi3el3Lm0tfI8ohOi1hrcoZFexNffoDyfywoOm+QeqS3hIDYO7/6mHNz24BfxJhjrxX
RYMxRJUToe/YPEEJfSMcRg7SWRSJbAv2mdnWCdiM/zBpxuFGGN0yJnMKwK7S0OT9AZ5G2FOzAzYi
iXTdYMCvwQduVPavf2hliKyhZQlRY0RYOtHW5GFzZxk8hIdC/IkeTIrniNTQcvAY0EQOMHF7cVA0
zSir8z2zAwNszp561s4d6Eq63PT6URUi1UDApxlJSb+ZP3vbTPA1WMIHcmou4nD8UElPXioMR3rt
dtyaK61Dmp8evXGa1YGNc2bH/ySX2jEmkaYvW49wvELQ85mNftYCaarrcOm15TULKR/NjS64AiA0
uQOStYhfvA4shNnI3qHuirq2dy9/0YyO0JPQ4tU4O0tpBtZrbcw9Sg/JRE3XqbyZhJNnXRBzlYFS
liu/c5k+l+PV+OjFaTi7Wid3wQqxWUpTa/EpE9rh2Rvfqu9m2LJBWgROiUXZKrVbYQ/ylSwVkozm
J3arQiX9NFiyJDhLpe4hUNUe1S3RVVl/DMJ34A3cz1HVnXWJ3xzSFen+bgpbzReh2jxu+sfPI3fT
Hjg6iXkonOwhOekHQu83ifqCBk6i5noDX8gwHJ7UMp7b5uoGNUL88HyTNky6FMe9y2Iz8FFkUQn2
5yBJkbSCj9l5ZH7qGoARqDG9JgJg2NXlv2iVPGRVPPrbSl/V4JYLHXXyeZO3RSXYuUNaYaAD3Dhg
Y2X963TEElnwUfhn3gHA9ggzAkEtow9Vinoi4Y9/2Viz2oW0xSm6i7mnH9dJQA50C/f/mWfp/acO
NIZhOmJPTaQ+6uvciedvuqdqyxhC+S27so9rF+i9yFBMcIOK85aDsYdlLEivkBKHBqqb9nBnZTOh
2zQ0ArclNSe4cOTk41OzcO6FsuPn5ltyfewezHCUCNx0Ii5LVZtkM9c0/UQbnAWjBT4x6GCHxxOb
2CKKh77I1mqTJKMYBL1tmFhxJuE6hRmo4G0uQ4oC3O9qZwqTqOb1W5hHNF6bdJx7xXSc2Ai/9Zkz
TUBa/TznqxdysrMaxvGmSx4kDGfPfelWh/Xxi4VqLqjTNTTVRXcvrnKeNTtcfhbGze8KZuGlM8Jq
u3/RdO3omLpxo4S4hBq1yXhAma/6FXFv6Ewv/yWImSzzPj0dGBRKtkNmpmGlBMQWj/bIkM66tgMw
D04bkCroCAIeMbONgKzo6R1+vQ8QP18Cj2UDb65pWubFOxPE/6AXnWeeUm04H+9/+T1pIpCV2euQ
1vHOAq8p+H1oNPRhbcCD2oXSyCEH2IkNz4e9f/Bsr08Gh5mk8Kwf6tgnXG8mIcJz/FilFI+o/2U5
lk+W9j/Phkf+0oY46qRmVhbEvShAJlTpUTuTmze2ZY100m9gV+0E1PtcLl9FHQOkioh1Bvfg7AbF
HhqS3FYTZGbMYlGwiPZ73muHwwgWx2mdAxm8BsbGwA9qX7I/crJL1Dw1047iEP1qMUDTgQY0C5jo
5QI9yzMubxt81PkFICZKkiYdm07wFxxsr/aupPQEoJT6uxFzdFZkOi+cNUZpaWmuMnmSSYlVOCBh
RRFosKYB0DiiQPXk8DSAJnKP4ijPhDgk+y93V/ILuRgQOqFmSXUyCnF1uj106BcYBMp6jk4DAPeo
SxDJRTW2wSgxSp+OHLITN7QqoqbGL4ED3os8u6+0s54K/C5fyu14rgjrNsNVbzACbnuRjtQHio6W
FOPnzRD6jl6Vaik3w9gSlQCBqvgneC+DtyKmYNsQTw4sWSmdt7oaNai3uNXUIeofPXZC71eRE+OT
mu51rXouPEHRlGNpfxjY4xlRNtZVkYyaoPl/poL/7McIsSjYE6cBFWugADnzEEMioW9gpvy1Ded0
vzdZgFiK2Yyjm3Lqf7AL5dIFOFjOcWaXK/MwfxJssM0KNajms7unw0l45h6PBQsexKZKFMPf+HTT
BloajqSz26j1Mb870+Wx1tL8OMw0GHkM+8aOqpZfKtHfBrhtm1xZi6YsnNwbYBlRlf4URX0+DwCW
l19tkig69IJZXGwt8JVljmmcYllDSNihi7jVXVKBYrXLQ7H8mj0sXTdfyYuHNPd644vtHROByPg5
AmBZIs3aR9V+YtvYXQcfkgsoz6RMB4vHh2SXRKEr46O6sPUeN96RiW3WBb/7Qo1CGZpadE87YyGo
oJL5LmXBWbJcYXv1NDqKt3E6P/NG4pqvUjCj0RAiSgokFYo2neNwRzd+XLnsOnE0p+TtLtSrnq4E
/r7nbBaGy4ax3zXqVc/evrQBz+6N3tBHDuay9YgcDoaHCPjT8+QnahtyLtNLVT+Cww/xI+esHfju
cCTvCImfxMnzB6AhyGR+5gkIiv0BC4kIMmiLLWQj13Tj9E+Fi3876mqAWa7aWkGgPO4B3vEmINEv
e6OjC1Nyko5r6nTI6IC0KxVJJv36lVmgWEpO+9M02m806pfN+K6WkCRMS0zHS0YfjcERlqucQMcq
QSDLVeRLMBRXjtnaJeFbiEjLSstlYsiFCMCSKOA1sNnJ3VXOd/EMJvDCJ++JLheBowyw3dloilXX
OKUcg+RPpSTXFPW3B4Fdva6NTGgbnV4mP+csMT2pcnc61FxraYt71yBPHV9ChNi8vGFRIkfcRFAA
QCl+5lpxLVo4IdQPtyHZbeQnlO3nh3lsxXwS0muzZYisnp6N+7adaFi5jd5x5uphcU5taEuSM2qk
p4WGW8bOt0YJ13twPnUt1HtIClptcn8JI1PiLo0Udq4yuLJJfRwnnZcCcGEUxY0xCiuIRa9lkDWp
NGF3wnO8obsq7PtxAHRElg9ARg9tXZm2oDiZ2Ucfnqk7AqbCinvHtMK4eDY7Dw5npyfnmriMVZ/E
IuJIUYGmcM75rDVj5Rq7oggmd/QIpkFacmloryz3k335Jg5PLLozLIQRZ7oH15s8vq3wczrHm0Qs
KEiJZP5AxMtptSlDBff6MdSb47O3Z7fG0Fq/bSB0lai3elXSX0kNfTCkbzjIpuOmIhUUWjXE2C5L
Ysx4JysAf6hfpPkj2utQ+avBW56yA38cf+H0g5nxCzlAjaQWEDV3jruYDeJV2jEMMCFvP1hjZ7L8
sKZddpfdAv9R+4MS6Ph4attpKFtw+n1gA1VG4lA6syb6iih7LlXOGUgklRXERlXTa0xUf+RbcRk+
OAzlyK2oT3Do6B7tX+sd1aQf68phngy/P8Ca7GUdGJv/Q4hyfgY6LMYBxWeqssGlEa+uZJ1+1IYi
qwqBsmaG4kGXonIvA7bPYWVbiRu6cBAGTvvhMRcEqPrJ0y5oSixO4+BG9kxoeOUYjM9420tat65F
nGlQDo/aqeRR5sFQHAz7mckCoprROvBZizVv8a2E2QMkL5zewFjHj6bujmeTfbhBqxjIi1Sv2Cg9
Zw+V8M+Ez7xkC2eh6njTAx1Yo8PnCVi5LzWiIseHyc05MT06eZHsKjlXOWAPUsPtr5PR73tilamK
hrMQv3X2sNzMaUzKzXKD/2yAXHsmtgH0Z63Vj0J5SjJQzG6iWIgEyfnO0ZG39zGzBUSuJLBNbEQl
9VvfaGQkYbV+Go1YnXiydu0r6UXvr0HXK7vyWecu3EchR/K4hObHQ25iv+pYesup7gnpRWgj9rlt
0sw5d0ER7JK62xGQ3iqVWgXxuWATBZ3iwblQiW4ZTDj0VRSRSDgaaUmlbJBZ0MuBlHe+mLlKO1Pq
sEl3dcXma02txvr4moxUgX4MeVtmi7roc3XZpIt9uL3Dopc+Dftto5DduP0+9m7Wulf9BMbkabJl
lx/N6aIOL7SGzDK7lu5QMwvKPu05eNQitnZZQsbq39FkQhNBENyNr2seEBT2ZSxAssDK1XE0jemZ
ZZQg5gdzFlme/Be3SPJfsvobAtQiiFpBppvhDMOItI2rEoaoQnbO+A6w8lYdiZR8+cZ1xyXGWHia
0m3yb423C8qbsBUrpbL3MjGVy3LyKv+VYCSnHsXvFc+1QtWLhaPYsJvPlh/dwLW5Oi9nlpaeelbH
x19xM63TUwWT8nb2ec3wBJQbqeTDTRFcgtE38S9HT06aobM1/Icygy15bD1UqXwt3JiMeN56Dwzy
r1OsrT2m+kYvijqd0OEGDcFdfjv5r2QmVAseGx9AhMNp88FDiTpS82cD76IfHYS82FVwlhwQZ7Tz
14N8+3bxDIOPQKAF51rkKCAhAyOID0vUTLdIXxZiQmLClCdvnz+EwBhlH46QcRtMYlikibDJJr7w
57X/n5YwLxVu6z2jgG8HAJKS8uFov+m9LAf+VcpT4i0cc6LAtR1fDM0zbDkqWVb3erwN09lfa2wP
sPA0+oxMj7O31vTaADgEG5mFicQZ41yGtWEjNfjlFM2scCfJ4pweh7uSpvM1AwAVs0yZcjRSSGeV
EYCkogKdsByWS4LsxCZHgNB+lJIaNQ/dw9ULPcsYA5sOdpsMd6yWMOH4X346VIIIkm4EgpQDmbXG
5TY6BUaI+brQseXw0Ny5LEhr/38g7fdgloXp0fYWkg0SWfIPrruI5tAn4LjKBoUKzGvgMygZ3iYc
H2dWA1AndleU34peVeK1sRUHPSFj+XaCHflCSBljujUIi3w0mc9VfzX5vX4Bt2h0wuMcBbx/q5pj
ETidasBIy7A6rY1/NGxKWn7Dti6imGE89O2x7CjK+aQsieJH7qSK+JKEbVUmUHMEGZudJiUAeS2w
/mzurg2Fck2wGDG+t3xd2TrDxxyK8TFGvtXdzG/DQ++D4BFAPiqQqCCi/9gE4KKbkE7QF1COzkWY
BU40+GeP3kKGdPinH38pJ2GC8C0QjH9Nga9y1ScZ+59HOgtWqm7sfDVQ9/IVZ3ACT2A8SV2Aunsp
ApJ8064ceGxdgipKZ6/w+wFS3GJKTFaeCBycsubpadth3dtn2NfR0buzgx6vpCkchXSrX2yWv8Dn
dYd5hNC6R1decJmq28FYhFcfRNSzJ+n7dli5vPTcYG66xpRYiRMMrOjx9pS4dz5RMjFH4SE9KgjL
NZ/3BHEAkT+xe0hc1mLui146vHW6G0epyCvm5hcik/qleELP+o1bDJ+Y+t11+AIeFyzPujiF8TkZ
2NdFZcN17xORZ+OR/sIS3F1RHsskLVODSSHefeNnntOhrpJAP29ISClzI2XavizovFD8hgfmXFs7
OXxnB3TV3IIRavaJceL7xmijge7PcfjZ9GIBuYrOP32JmO+6d/rgJBA4p41nkfyPbdOvm3EoHov7
3CpPgX7arx3yGBJaJxQhxww2kmeFsIZ/zAgqddEv2hE7D4FturH2cip/VSVAJtIcL92xk+/2KkG8
UMhQsThvA+VlAn25ELCEMXuMV0OenEtTuoCVi1qAe/sPcxWGok2pKgEUlue/l2GvDxp8QEVSWKU0
AyscsOldfQpjQg5hMdoqKAI1KTlREwLcFBx3kpRjF19WwWLsqSkF97fBuZyVLhupnOD06hqbZP61
DOL7HSJjEj6TRfsd/vFmSe9yrQK7JlBfBnFzcmbS6CbEeTe+TkGtGg7heCBbzsMSj1AmyaFCdYkV
gPxDIF7B+oODIKt3HPvViQkIiaOezQYBK7quYcXYadnqrI0HjB44lSTADw6gDylKJEqzGNeqW+DJ
Ob5GF5liY+kOBKKtD9dDCRDI+56nl3ZV/H+WvpTK4sKo5zZQ2vHy4+dlIBB4ZPsVap2/1HFRR3w2
7GvpiCNSF6BRmpTFAvuqpa1v3/iqN6upmwTPfMaCJhG6Jw6bc86Qa7qBu8IJh12+zmhSjjhK527F
dpGv+kFIxXDVqTnZz+csK8xW9g9jcuy0EsPdTIi/9XMFV9OzNtEsH6tXLF4ObCH+n/tWdXNHz46f
hpSv5XaEqhOrdkC3GQAHUOsE8oFGRXEZ/lHFy2rfK0Ik6JD69Dwr+fDBcCrcFZwn3/jMmcfj/V8L
lAuXzLP+0Zl9f5hzCqPEvdU6zeIxlatSsvtERZq1tL+9AG916DudRmL1Ux6T6b3ZKGg6BE31dFVI
6VJHMteDJHMJNRsFQoLdTCLAmQmFFcA7/I0qGRLtBV097Y7GpXnGbp0WOEsTM25yy52AAw5wT25g
i8lcdD8zEpFJWCYPtM0j9MtZgorwI8Loh+ldLiXbDGnYMLHfQZdMhfNDDK2D86waXGh+V+HoxrxF
qAYF79M2ye/xijsuWSpZw6xtMo32TPTd5oMIspgF6e8FzKqXK5Vxn26y3C5c24MPZCSUIo2v6Iaa
mjC7qIDAQl9JK/wDDYswZYHp0l+Uq73xEt5Q0PsOJSAwN1+3rwZv0OqfvHUqhSWg0Hn0wp9hrG61
BNhGWVK7CdUiHis1VDjbnTxbYTf/nmKWo8g2GQ9nG8mpbRwG4At+lALX5jxG0+gYK2xcbD/Lv23E
p2QyyeyvOrNAc6C/yW3mWXCGrzPGyTtFJHjAvaYOLtcb1PNSIwKO845EVvRm/fESy0JKOUxIuopo
oHV/BkqMJ2MJw1gorL/7tf6vvv63W/k2eGGjqWCmGKDUUVn4O6hzOulXytCqOlNDuDzL9Jv9zqhg
LiJETmJHdIPRWJE2KGRaSBBZCbVFF9fS2fSUnz9RYhr2GPkYiH5T3Xs4Ll64tn1Mg0eZ1a5TsMAn
QDgc5h/kQ6yjXlqy2tPND7acLd90S0mJ+yAHyvgUUH4uwgdR5N1+dHeXRmuMu2JcMK4nSSjZeZWt
hOz6NIQCSk3TzDrTgTuVNkeEaVvjzk7HdWgiDRAY6d9hCT+UvScPcXZT2BoqWDE2J0Y/YxwkdYXF
xJ8D6QpkirUaVGzGb3w/7/UdAw7+tgdrVWXFqhR1S+EkQfkOLYmUfjKnU8D/v18N70qzEbmNLDQi
nrsSaLA4GrmXGwKFfyeRT/LgDtE4afJ3I5aFqUqS0jICJTjMxYH3sXYcA41xMq6aSIPl7yiz/KfZ
pzZqjRzg0AK9d0pQ5TFqeCsQutvUWSbGFtTlVDLvu6S4eZGTdqfSvclq3U9L0o6GVwKo+6L0g5ZU
j1UvnZb+KMkQpuhHSbasKbFM+hTV7TN2xgOx1HM9cn62E8qUb2nfOG0d1gmMyJl4AhMzO87Q7Msv
jQTVp0CO2ZFgiN+ygDR/YjAZfJMpst53ZtwiapO0qHdALtUuyYiPEYgjcNU6dnj2AIpNwM+7Vsoj
req5ErBR95eMZndFgl4l9DEoGSIDvynAuEVWvw9fyeVaovnQNCbVs4/6C2+H562e/m7KKv28N6Ue
nHKo8mTmVevjGrcDYFjm0bmK8Ai1cjekkd9FR5K76+rkF3FqfyzCtd1MIbiI7JSUh6ctjeBCIfJd
xo6S/GXGI9RHCXV2pvFf3EchZwBI5B0Y7QaYi1Z9qAXiQPNnmLQYEIIim0Yf18M5suBoRtIBjojs
udD/vp28Q/HhAtCt3RGpigHXnjIkPfSfJvApTNQFpsvfl7QgsmrEt27J4AS2nfqzde7chV/kCwZ6
ai4v0CJdo8C9OIVSypiLEpjHLUVkp0jdUlJBP6/Qpx2TQDF+GZEYAxOArNECJrftLVyt5wvOVAWF
UBli2Tr/AAQmsqGn0c0uvD6bOQHqFA3FVDdGc6QrXDCFkxX+58yq+VtpZ+zyygG9meY4WuHYiWPY
YH9FpCD8+nDFnzvrQpc+2FV6jEKQ3qOCYdLYWhVtA9rbQwiFsQ32JKddM8DQ0XphJWUup5mUfyZy
v9x9Ph4JwScOZ0qwG66SvHim8QZYxz8mEdpxz6CZNCFxghoIIpLqOMzGBO04Sn9Dryk0EgAu8PJg
ZTcPhbrClewEUk4vlz8XyQgygtNQ0V91L1Yk6Vi/6MKhKFdP/S3fcSqRkKk6Ly5OZgGQeWwGZ+St
0o0cKhq8uox4XvcyzRYbku3fZBovshAQQI+QY6Z8RBSmSDZPii/A/GL5Wiy70nTsN1MPtdjr4cVm
r7yoWJnTrfgRQQU2AVmCfYTMZBezs5x8+E1FCcLACKYeDPSaXRIQjYrGDjJ+xshCK8YsxvW0BY2u
Ldu2O0HV2Cc/FDBPD9iDcPHEZBX7HqKxPv1akBvYRkC+Pw8X0nyiTQZrOQjkCIggUnedgmRNQfwU
WJrg02b+6nPiJY3V2BnPBR3yV1vHAxEFdwCh57lXfBqrQNblmh5TAbNkviiaWoL10Oe8rBG+T6QB
fJV4kPaO9fVscNkU0x3KL6oiB6RlNi2JZyEGgdg1l5ZJRaT6Wf0OHO0Xg8gYLD2uHTtJ/VTCgiC0
Tr/QyJKgIEJfCxyozo7C1ZNNbNMPvSFm2V5ERvkrLOUiTEexbUrBPDzY4+S1zPrYkbkbzRqJto6R
hcaP6fa4JhEXVogD0ooT6wYE2CWH/lYnk/JWrNAolsa2JPmB3RMGQB1VbGsLUatg63y5QYpjIjJ/
nI79XB5YatbAAI0mqnWisYsVRAt2c3yioqQjRlA+yAnlJaOdOFLSVZ3mB7rkLSkpi8eTAMo3PGSf
ljpEuXCwE7TT23TWnQ8V1nvy0GJX8XnibTyMo2IFmiWE7x0KFmnd+1ybVOeNLDcvXq8EgUrwMWsa
XVf6HbpgP2QnHl8txHXpWFaEbP2KWr6e3ixFE8CrrAFIqd8pI5Z/UBLcH/OVSKm1Am01raisA3y9
Aj90XFvUG+uwMvcdoywSn1HgcrVJEfxRkFqS180kKRV7ESPxI50WNQ8Kx3mO8cinaklV+Li13AFW
fVCRbBSKVz2jOCz+jKTVtCtagybnoSG7Y6Kbv6bYlrfi+1V+sQfVemH371xUZei/7cyLHAoa82Fn
G639Kh+Zcgw+0d6oYXbLTSHLDi5jcOYiDF3h/buSd3gdHghrahvLbZ4XdvHEXs6jfoBosSOfuXUB
WEHvxrSHt8M/ObUNldcZFHimnwz4eWdkpr+gIIaU2kebEE0L7tzz1ovm6S9UjjEgNSpMkWWrjC1c
l5+GzsSVz9XyCkYFVdr4eDNMeha7JVxXMtdSDqDtHgzEBZYRzHO3hkTimpTCnxydZ4xSk/gfRAs8
ZlRyc5mu0CG2TJWD6IKXrv8SsLz2k/ZPZr88S8pscDP9vdn8mzGc2L6msEV7gsKfgcRV0KLckNWN
FuAm8zYSYOQhr+Ejwn7OkXh950DqYALcvM/tOL3AbvSkZhNCtWpVtePzX57TFtnp2/MVlsCPomae
ZroqsFRbTiA5zKaoMPHDbyTGHuBUjHKHz8a2Q3Cs3G8x1bUvcx/o3JXjJERUsH6SBtQTnkmhK7CY
0I2wX2IF9Lww1InfdVLQ7CAPIVq4kDKECGAd+2mwDYqnmmIu/rPBLWy5voK4sBNRkITkbUX0q04B
1UrpL8NC5g7YJTxVuyfRFi4dKRNqE03M3mQNcFIpJthelmZyEL8gAmlmbDhJ4mWeTedIy4GYe3U3
Twc6E59NLZSkND+cyGhgl5V9YYGjeqAsdka7ESxYohNAP7gL9I7xttRr5T0vxamhEHiGVDQXtNGf
ADhVa4Yg1+A9sM+w4jTQplA1vaW2soqRkJA8vJxXzxzMVX9KtM9I2ut7AgiBKchh42/qbQSfGmAe
hLKlH9mx7MeOY5mxPLxrAcUc9NsJUlAMXHCPIExA03/hb/MaChYhjH+NMgT1krF2d21OtmLR8ach
Eh2b3fPUSFEAvQMnvmUFvU2isjbEdy3Ub6gcL1xenIQHE0D7YdFfQNBSyGCBHURPCM/kI5OsG1TZ
IZ0WBaUq4zyumRKCa1Df0ThZ90oa5Wz8bQckqXCFBAEKaofGRk9n+upA/MfBiZukbnLRJotSEkIO
MrZmAk/X+AGMBAqVIZlwnM/3GLhvKA5rr6hGkDdvxyd5/0xcwarHkryLFgZSQ/7oL8+aD0sWrCdr
hNtsxS1PKjXB16u0OOE6spDQiJ2iSFlINi1FSDQmBqlLBSIw5cgiOBf4mYzSUX+8k1gkNKcwNE9B
fpVIQAM0mYkzKfvHWxc5H/+MdZDEECgojyh6WH3pOBI8029x5oCpPYxWEDB2u38BpEm0WYRUzxLY
qmK2rnAAuqnUelQCN00S0pT5OCV3v+LEZBUCrv7fpHEi5bImxuV+ObbmGNUG2nBUZbmIksANpInE
veDpu2wcb1jxptToWNpPJ4vPGB5jSYglFUBZ77XB74G0qXl67+WEH7u56w1HaVWMzse0nS4W+CKH
b9u/+xafA2dl1LTGartKcMmN7zzdR2NfWverEvw1cGox9EA0isl6t0djYFeCbshwyI/NxoGwQf5t
TlcTkoQesf28BFGqX+FVTsSKdvfklPKQJBq/NaI4kmhP/83YBJB7jFwA3RmMoRslpu5DbhIaWcxU
MuOzkogghdJOykvJx3MneU7VTjsNFKXs0YlQIGJzwclrUld9McRbwS+ggNfyx/GKfVKfJslZGD0a
G7iftzbkf7hGqZD5/xkUEXVKu4FyYDMlBnjJYX/HeAprAHuqfu3fIF/Fl++nRLqOGwbZzs+8cOfU
SrD6ut70K1LF9jZUVPbVg++RxJ6FsQEjkEA03Y1w/ULNTwStMeUWpPqICqnq4swi+Hh7NJUAQB5l
zmUCFb/SxQc5Mjnlxmp0b8wY9p0FakMhkJaIClkGb+Wl0SmyOt3enGchHWnYa6LqQohhYlCVJn5N
OPFcLAlaxyCclDm+V6JWHd0fOFaARUXAlbeubariy67hWNJMyNGx7TqAsJAPSR8wS59zLYuxY6+i
RxjpHWnoFfPALzhqSH/9YMw5nCHysgjodcJ4LHEBxdKfVOoBMwT2NI8CwPSOIeP6YUXDekzQ7/uR
nACJDdJqibT1rNLWSR/U1FlbpzQy2CzOJ8MrlvBlC1vQfTYb1czsFxm9JYGEJhavEFwkyk1WxPM2
tgRBeSHmWZ1SOxQMu+azOxtA/dgG65AYwJmrPzUY2vI6v6UajMy6zjQR/Cbda+JlcKqWSqd7XhWI
+yRn/eyN2joM9MlhfsXta1nimOQmvVms+ZAGWLTKcEY7q4mP3QMvlqGYkaSxu914GGyFh0I+kxLZ
2f5GTHQJp5674zc4dQ5KzJDHFGmqbi0uzYsudc7m14RAaJHnLT5lcAZuZanV4F6FEIIqxmLuorm7
Cr2yi+smVrwT01tSbxkxGBBomC3RMlTMNlRIDfhJegnMCfu4PEm9ggCMQgI6u8Ca1qZKRoNNulOj
3zo5EEvm+QDUSUmPLxehPAnJSR2byRBpCNlQ0303ZLWwgU8RutL7TU19VhgGTtAK1ojcbXWGyhHd
7JT2RIoYCGLWoJPQ/JgUmjJ/1ou1SdarUfGKxGGwPdm5Yhvn+WAquyy7tn0vbV2VoGH0Wmmz6D49
qo1n0ukcGp+USemHB/cuTfTIOfgmz7CDby59kOjbrfIgUXB/O/BDuZ469IeHeq1W+4Z7ugz9J+Jj
wstYc656kA3/7O41K3+Gp/j1+pVyQ/DGRnHzYt3f7UdgDXSocgeiXJbJVe9xARbtTwyqHeOhxaaO
vM0TtBga2pqlOemdfL9LGacc1vPiNfK/BQSLKvfkmialYaA85/Ln7Wvu6AxecqKBS1M/9hAfIeBm
ecLwa5etyjMsFfLIV3no7Ha1Grr09TOp5OEeO8Z5QmelHWKqmad7fzK8UXv1m2M4hvPDv/r1QX2U
2t8JALZwEzL0wSNw0ioFDIKcynbI+Mty3Lzw33jZiloMJsPWoETmUHm3fhJrVPXCdtAKtBplazu5
MpyHxums8dlu7ZKE+HHKdTNEOF4POjsGleIYWHFLTKEEUaL+5s97Tb3siMMWEPyHsp4K9d9/flX9
YX1hX6mVGcmoU1wGZBlNiSxM9CeazM+HJ9RFM3foV1fI4vvjEW2q/8AFvEKfwUPZBQ4eiXuspB6C
dzlhwy2t7jnPXk9UBDPteoTnspQWSl6I5DPl+2WcHN2d41sUmFeDYF0hp/8BMaHTE4XuFCSwxdN2
dVXSgyZZaieoQsgkIgknMwbw6MF8SbygdnC//XJrjj0sSYbEScINtbpcLB/kiwjKC8kFhR6aJgG8
s3ohsUKmhPye5eZYV5OA/oVN4Bz2WlgSz9P+G8igAbf+jkKzDQMB7g7nSn9EnAS9ZjSLdqWi5hjc
ZBCh4pu4sSi6dCZX54Ml1GrbvtupdcVeW1kUqW6rLRJcd6Hps33NF58y+ztMu4GHY4+9tnkmKOYC
/WCBFG6FdOVgyP1AiWSyaMyZtPSxDwvdq9QRvmM/NsGtRYNxPj75veGBb/7HvwBW4rq5t2P80Oau
/IenRa6KlvD/y0LXJxuce1hU6JgEDnDY5cLIVOoDTmydA10zuuEJGbmt5/qt7BX0VyxidLuYeRdG
QhRBHtXAtnb7JGERfAq5/STsmN1N9qL5mtlpD0ZHfDP0y3ZB7dW3NvEwzL9nKSQKAAffDzi7IkSx
+KS9j8LqApdRFYg8PvQ6zPN9xkS66UhL+hzN4utV/TZ1FJjIzz0Dpo24l9E8FYzSjfkdfxQeSFsq
GSRbnYOgu9aiq8AZpCFNuNX2LZo8TEMYX8el/ygI+uBqlKAS/t7sQmTVth51Cw36EySEh1RmuEXi
EaNgwKAvoI6b1ji7chbBXPjF9zxRV3t8dGSMDlykT4L4m80SCjWbIPtX6ktblMTV1FgR754HrNYv
ZsIWx9A5GeuyO/v6uQWut38wNNxmFjefrHb+iJakD85U4iiyKc2pkoQVZgeJhGtxNsCrqfU8VJLy
2OBrFfsiNGPlx85kaIH0Z693i6b+Jga5fPdBE8FCAdwdLbbqmGg3VVcyGbhLXLtzRM9OFZX173aX
pQ88i0EymvVC8iLNCKoafF/JXxqKPakg2K3Mic2DlA6feiMEED2PrGKH9cKxjBzmBrCvnI7kScXd
VKPjDfo4tNHPkXvst0evGBBiYdww5v7sMt8Fe6xjgKxHZWzzBy9/gP587jZn6cv4kIdODSrcBIwA
OJ1LKGR6tnD5aBDPgjxBcNKKUE3zdJkwRPD9B0iXTUqPI3qPnLYfs4nlteEg4M4LdoKWROUVkq/H
BK9jXW48EtMfCGBfA1r2dKeWsYtPMD0VBmCVBg27cSLBGpDDW01uCjgmct9JwcZVXfb6ShDOH/ZY
3Ud+jMNTvWMNZXic3q8depFi5Mh9/YUqqZfp1Xca0W1eSvHjGMDBepmClaHMUQ3tYLVpRtk4hxlH
R3aZUqtNwDETc9wj61+YqWq9u86D3VO62A2mMuFjcydVe/AImQG9s+SsAZYLosTUoOjM2fpyWhiY
VG8iumwbFsvmX6EwRGkBISqXfoUlfa5RD8rYLnXQaUk+J+1yCdei8u02wV6egjPkmgs+YCilp0Df
ZR5E01AdWPPTWcF1f4+RnQKZGqQ+8hSl9MMZgIfJGOXGxE8szHee6RWN0m+rdBAY8MT9EP1uEK80
0DOXoVWVpNZIIF90DlzynADeMajkWpIEdldBd85YHzT2kK4EpyAo6vLDvWKaFUHqhppQyKYal8H1
3zUg/HH/cw7JQo60I8R5o4BUm60RCQ/e80x6M89m2wzA/SleUuEfTRD8Eha5DY82M+pkoYveAK9E
NAhA0Qv3zroxg1sPXDyrNxOs/gE0w/xDp3cYkH+VUK4R5sJA6QcjC2pTSm7VZb2GY91fvPMgXCZF
sm/CNEhgKoPgARlFpCwkwlzrDQxS6Nz4/dKVLPfbrADtOKjvNJ/L5L7CS5oM23TlESKRA+zw9rWB
a+xvsMKkl121z3Uy3TD0WnOMv8Bj+/KpQlkzXMJ+xCityMS6TScLkxc3+CXm9HrHRtBrxD2o94gG
8oqa9QmH2a7R249Lp+eF+LjoOoVkF3D9b+ggvfh8Z4rxMWBJma3jTO8kNKt/OUnJ56QixnZ+sI3I
Mmpwzca1Nj7NS4VJO8bo60lkn9NzSQP7rZ2Rf4feybf0FEXegYu6RdEiYPS/jCrE71CoM1mT0k7J
UCcZzqAWqQi7ycj/zXwzdzQM3NtbQRu1J1FWMddyizfxrVipVzhNZL6mKP6ar+G6dZmDx6Zb4y9u
YmsPy7351aTKUjLyHHm6yhdMroNj5wfllSvL5Ft286tLDzYXii21tY/OfvvXjjuW7rHftZPylg1y
otb3hcsYL8wFQUKNe4uyezLJB4n2v4lkj+5vkOjqOpSkdT9sdmCnm2nKcgk9NKTxnlmMGF1nXxdm
8Q1Yc9jfHowVWXVRCAMBMkV3i01TO/RIAgDHlJFwWbW3nAN8vv9hqLjTC85H34zW+IxbMcI4XCer
Z8tuSmpOe4ofde7rb8Cm68mH4mcrdMFwfx8ag6bznmlQLHJ8EXhpTbdHOBJTv43yyuqHSTPPHRBG
7PxjlKYx2CoJQ/xkIFA+M1rCsaxYcPUK/udTGcHzDvTmtpISNquBsJKn3YhiqjrXCMyiSP/dR02C
wTnbzd/4YEot5KieHIn07spb91zmduUfboNC0tabUiJR6JWhxbfFVnkPrVBpW8Xi5cJadj/LkLl6
yfrstQn92aI0ArR31VvVqlNwvKFhdKX4RSucIaBoTKP/k+4AewVmIi8qwAXfIIKy0YvQ5PmPjIPP
G3/hhtV0kqMPWheYLZcUVtHzgKLaL+osp4Njb+hMPG/Y+PxrKKFEdU84KpP5MWIHkTVl+I1WplA7
4Ds2u3Ph07wfcrgfh0sIVUcWy1cfefLdAGhxWiVpyi88MoPuiCpegsKDz6VrJhWyaYbys8+Mfn9K
XN0miSrynedzeSnedGeFRMWnqi8DYMVTV/hOm5V+Nl1L4DopmqxOnfqzGqlHJn6PTDBL7ypZEB6k
hpqaCCU2coDLInE8hvEXwgg7P+k4neE2HUsxM2sRE27DwDBiO65Jli5zmGJgs4naLs66rt2XsqmE
uD3fLyXyd4lPoO0c4lMA+d3sikgJKoHZ7x30KKv2vAPbkz69b6wfIrx+8XuGFwZ8JKO62SFguR1s
Q7iNQhwwuK9JwAkDQmOYJ/4Nn46f/fo4Z8wVLWoaaxbmzKQTvJ5oDotIRvcd4bv1XV/CdIUh+1Fn
vmQhjDOo0V2xNf7bZ0mVrDBk7bpplFeye2CN8tqtXvJLNEQHlchz+DtUmC2V7XDASx3xadKai8Lo
Plvge1XoZzp70+utCXvbfjBZDGyRu+NTrz5oRs4U7BVPfx7V1YQ6UqSS94B6bk3U/yrAjHoF7zXZ
bTZinmd5jLp4va18BqI4HcmDtaYJliP3Gn2TOrUy9EXhJWAXHQpy63MIn6TmUyXBtLVbAFVOS5DO
V1igxDA6zuUHrNg9HZ1x7lljBXYobvFLXEasrmoJlZdxQp1uzuVR5WHd2fM50PvbkYx6q/GP88T8
U7KcaBnTfkLBb49NFkwE358O8QH/GAJ7PUinEwuNwx1RJvZNZgfhFWirVwykHCCu5lMTxlzr8SO6
H4MtRqVc5Meu2hpWmG/CHJrbNVyeAQaxZEfCiKyDOcHbGPJcg/IgTsnGAeD1+i4HwJ3LKkB7Z8HF
8M9FsuVoL5xHUJgiMT0wvq0BuNDVw2oZN5PTlBaxC8Hkd4UBkZ41KhTaVdD7HHRrCFv0ud9FLFyX
vBNVAoV8ubxStEc/pfMnA3p1Ygj1aiNWOgqidBiYeg7bdnPfb9+G7lPBBpDDlbL1AhUXMVZGHFOG
5m+zhNcaIK7aX6+vbpYTYJ/pteICQsWcH8+5vcteBWPaZV/tVDX6HEakD3EPUsmfHhw4a1bVHKOk
H22xrU5HYeF3JuBoW0pL1i4ZLBSrONU3foCTPV53BurQGiveRICPLb+5JZLCtguTfccp3XJTVP4c
o+6INUaGvY/Lu/VV89XSQzXUjlqKidRCXLaJLcEPoPZmiIvvYVGV2UMOsSvOjMMSOIeri6dOipFh
0hsh4zhEWP0411HbFpYs+50x/5adswz1J2vP9siyB6DABzcmdfY/9mow71xNcNxtx/MFf3qWFuHC
YNesQiqlTU0I9YnfkKt35NPuelmPEvfa7jb3rvpqs4Vs1YTk8Xl2/aGdIa2tzqxWJ9Tv2cXNJAKB
eEN6jnEASGtoaS2MzuQk4BUSQN23R0xeeMya49K+sAQ+VpNWKNk4+0mlVLUaXMgy05w3Y6IAiDDa
D8iAivdwQMpGaPuJHtHADbgiknHz/2RvBYzFAi8qqDXbTqk54qTCWbl1an+L2tNy0fugNpnvZDyF
A0O50Bc4GBLPfYuo1IGxyPYcHb9fp37tkjbnS83IqK6hOAv2C4cvBxYPAhB/7jBAZ1jkn7vMR2oV
uZak+ry01hMdjY78TZfZX2dXWQBiK0U5n7t0eDtWC6L4wnQGrjL+llwHcYkKi/ZVqT+Cfxk/De1P
jIY50ud8RNL5Y536BMFG6KJEG58sQNhMmr/5SJDhAhrTMWXAMRVc2JXqSwXPu2EkV8nLLHrp4ceP
XWUj1ZOeUtpPV9lUc6UY8RnMM5J3hcscAaSNqwweF9h8RgrezztYvEYnB1gL5nGjkq4EweeGXHNc
YDTFWhmCygnYFOBpK3E4BQ5p2C0d0A2v6MDSgkogXXmgiwa/Uhb9PR312t2MenZzJv1pYGSp8ZGy
AhmVAzUq/42P1YvJ5Sicy+PTXms0iQIrqlUTEwxXpRTWaPS3ipGff+FaMEUHawWab40rFxxOqr5O
JW9Dbvt4wacNbe8IeGW20IsgEivH22Ye9gbj+R8+vrfF7VGpAE9XBa8m9Z/DnaCFveZjDQSrREom
vx/endOIT+XpKxNcNXihcn6lCB9GOHCC6Kw3VvnK1IlGP1oLAPvNYiagdgD+s9VtYM4NGcSgHAyl
/nJUrvz5QkyNSeDzWBshGP86kzRwR2U3C1xifyuYmlgXU4+0/l9nGwImRjogl/sVYCPl5xhI/qXQ
JfB7H2OQBp8cUdQsHtl1NB/yYwHjHqtbTc157oyVE57r1KrVtD8ZqaUt56ZuLelWh1q+JL4racnK
5UGQBXqBMy98oWnqi8GTgBtefp8xcpoVpARrFB2E8mEhA8VLeSQDVc5EhfD279Sj4eIMB5ZFjvSP
DelRhnRaVAg+kaS3A7vv3wQ0oWX7I2EBw9QCUDuUG9o6V5tfFJ0kWDd6eE/5RJyYvLLkvXsWLBV4
0Ixzx5NAdVUWqrfX2sG0h6GJJ4BEyWTh2WG3wRHMgIfur8fs+w7qULsc06knhYO3MkIpteSjcdtL
vu994HR8rXtw+78jDO/9LAD1ka97HsDj5kxmCQR+rttkoMSJHacJrxVgmp4aIGVA9n1ZNV2ogSy2
hj8TXHFt4PnRJMGFuNo2LhhPTdVT9AYUJdYDk62tm8ufZaluxCj/L0iLuENw2Ux2+JQQKZBJzgrv
8YX3htB8j0SPK/WUTAkAbMaQ6CSYhuLtHC7Sxd6cfDajs3cXuH5UG+h5vp4OASMp3rfUo++lXODy
A/Xmhjt0IwPlY+nv5LWJcWsXrGp1hyV6QS3FfRKoEy8/zWIOjV7A9PcTJW0XAEQwAfTHq1Qc3MKE
J1CKLEomQe//O4ab245pt37RiJDabo6wRs7AT8g7SG8UbdKXxLR6Iwp/ZmbnSsnriMfPLwN5zWQX
4bsW2sm0+MO3Dl76B5GGhWMNxWuobaLXBBb1DbNINL316q7M61M/NgUY5YNuKFajTsxQtbntqT8G
fOzE22kSVdevsm1YPxrdIX6j5U7d0eFwQu4bWu0i/URLIf3nGxrqpxEfji0TnobgAe0B7ihoGptu
QJN5qXJNie8fy6UfV5RdVf/RucKXfNyT0fI2ZPl514Zcabd/Nsj1pvpWrHc1VJRNvrDloscNhn/U
d8jF4leN2P11PtAOO4Bh1bhjWu0Qp2d/DGc7oofkbLY2K1QkfRCmBMZQB6tzCi8sPP2nPxSHb/WQ
r7Wzcr1WrsbHDEfGkvIFYVSGkT0XjFTsVEW4gnLlo2RNH8evH0eLO8J56IkVycUriGp5ss9BSM72
vmJJstgqHujZnxrL0d6Qs+84Y/1cjmNSm9br3vxFAYtdZQPaTGQlSRtCOorHhOnICRrwie5Pi2R1
89zz7N++oRAbbgtW+MNuUnjHL60hLPS/HcjY0Ipt07MX7QnBn03W9ltZ8FvmDqIG9zWd10GyPMnr
da11Cuyc5VZkVQU5unDDPivgonkA7pueZ5Jt9eFE1ryJS6C4o4dHTL6KvdHAbj0x2UEZZDZYiEu3
bAFn+ebkgkwOzPXMWD4rtB/KhgO2/+s9d1XIgGCh/07tLUzfEXMen5lDm8/Yj5df+1CMtv9G02vt
ooiotliD+lnvDwT1hkOlv95u0v0BfdwkqUdVxgUPFo0iSiHslyTp7FrdPniyxMkY1Mfvj2Azu2F9
Xc68ktC91jbrFdQFEMDuRcEvvsTkNxkjHueLSDCfUSJZWoKrAYwMVuyPEBTVzgCeqRQkgSvhqA/3
pXpeQcF3loqUvHQLmJP75IT6kudvulgB++ITUUOsMqSNgQIr9QMdgKQZYIwq19aoOBA6v9TJB+iB
LsMwtdTJdUxWHUtBBqZrhCzz8ElOkgUi0I2AaZHMRNjjVF06q5V3Xcs1HtKbdgzBxpHrdi36jcMA
xtYWftgHDePljVfr3i/XneJz8DIwwfK9jKFP7l1zF1c+bXK2yIwysyKFI1MxYi+K2wxulyekJQV2
9eTn8VBiGLfOk2UA27egyIGerGvyi7/DXzj3FaDPa75lFcTiMUdXckoKhv2wjVedSOGjRNGGk3Oc
6nhDEOSHkpkGOBG0EV52P0ykngoi7TMhUqFlppNeE2OqHbca/ii63A2FETLoxcTSh+bWyMXi7trb
7lO5rmRhQ17L4w3wzP87Z8j5d4lu9tYz7PpvEX31Ztoa14n3uPQDjAW6Po+wOM1n0orMOeP67hWj
N+OKky0T08oSuK/l5ub4VSIbaJa+Ybg1819D/jdfNl6Yx1NFGE/AUhMjguvUrxfRJb44cVu6lWyC
PmZY6CaMch1+3l5Rw960V/vQoSs/7qhqhpNg5rsOtH0Yo6QjDwOwh6k85HX2Ex8vQjQ1tgb/8z3s
TniUlzaDj8y10ALy0SdTeb6yZf490xL/xysWyzVefqmE/kltsStsF6YIfJPLB1t8JtTT43fy3SR7
k2smiUX1XU0WTvLoJTkM9ah1vlt1nGLBM2/P11w3bLp047VnEYH5EZjXyod6rTySmahk/jsAqVam
EnICp4LTX2cB2N86gi3KTWkP+O793WgrtlYik7nO9t4+QFpyfYNF2wRxLpV6vDhGOEiG16WUgbch
7JedN1mXdz0THRlYqFa1kMgSPnOYkVDy3Cxc2CBkhqk+K5PPrJ2fCOyB5ujauPl6h02BSUkqzNmu
tB9Ou86sEGYBKxszgy8lfPfYupESuMReym1PIPl29Xnj7uGGoWrnBcLpmIYUJIqxazGua5BS4+4l
l3iMy5mxS6YBxWuOumhmT851pkGE4zRRVyXMd+p8qVTeRAgZMMmcxMEy0rNdk3xacwO0IVIqxG92
FmEDDAoUugy3RNc3D7a/M/Hl+8yJxJ951og1TG+mSVUG/Klco8VPELpD/A2HF0McxW6oSw6mdJRu
K/CT5hgVSybi59PFnR1AVtPNDnM73eEi7qbIXICljPxPobXOerOCBq7qKSsJsV9MbgU4uNmGaEhl
Ujsft5/TWFKW4MyfaKws7RpAaLa5jqKWSoJaU6n826yp1dzTh9dxz29rPwGbH9OKOyr87mq7khCn
mn/f+9Yba3mdsRvuqDrt+/UsKbJigMJ/Se9k7DNh5W3VT/MxNQsmFAihom9meHmXOScIXcq3X1O8
ZimmqtBrIySeW8VCyVbk6MI21t9g5rRUp3NCQ2ufChetHeyWQO51D0OaoIudNd40LzyNW5Dtzw7r
4eRfTkOKW92xBzFgvelIcuTI9nZvaBF51749duknbWPMNMcOQe4kR4GCBhh2KH47ON0T7m1S7Pxq
oyCygYwEsyWcvIqYsO8WbnKwmOWvv4rA8UVQFjrCgEwfZQCFwY/p8KirmDVSyZiVv1XVCqeZL3Yb
BT6PKaJwJmjJXm3nXvg088V1yw2wD9NGztuSP7ryVKm2dq58uwn6d1hCcoNKdg6juIsdzIfzgaUS
kLwot19GITP4pHokvQG+J6JoeTzWxurktUZBo3QzBLL/ZtcBBXvBm3GkcTZ/nWeUXYPbPQjP32v1
68EZPOVwbq+Yb3NmQXPp8jnByynmfj4xpjITKY8pKjrDdxAeoBs/iFbkfzKjxCTB524MTS/sWNZ+
B1UUwUf/kTnGjlQT02rVhNpOl8DqlRNixETwTv//BrND0tVvxWmOVlpt5AjJ8DWsmehEhT0+oDDL
48bEsRtrV/KW6GoYTjsVsnSw6zBtISOFzG1T4N0zZUesjy5swViH7YXzvKBGJfh06652nknoexYx
SuTAWFwBllOKf2qdI9jgnjJEFUK0TWfb/di3KU6GZMPwAsiPhGWZDeCF9NcKGx35Mw+J279ryaxV
Vu2Qt//QlMZorQYyOkWDrhYic3IykPRaDNQKqsYUXFJI+jCqTJpknvDTpwJ2KU0DgvUMpozVTUee
S8/odC8YgYQktRpge7sAmi4ssn0a+mlOzNILBcwCQVgE3jN/iierO9QEM3qbO6RAT9e4+w+GEp0K
Hi/A1R2BLVan0Hl2Vm1jQE6O7ZpxSk0K61/9SX0QjNLZgjIUGmsxrMMwxRW0LkIjdbML2OAu5i2A
F2SI2jnZR4XPwllAfFEXcseOFfe1lRZ32ZSSSTCW04yFaU3JdqR/8nb6rjeTwkN381BuNK88Fl7i
feBqU3golvsraBHi00Jn9HuAEd7P3c+tmWigZwGnWObP37AksWWlnlq+Wy0wWzHjbYOzwiEUiY/X
cZQ87ZJKNfawSpx6i7dpYU9ySBvoze8q6DggzaqjBFjr/bBjct7lM3Hv+SMWm8yo9gEqf4nsoNem
ZLgpQRoNXIPFQfuFSX/rlaX/NDfZjzDY1yJAhUSgiXytUOIg28yneAiEo+0m3pvMXColHDZksgFk
F5WzNHRAv0txaVny9n/2V5kUkfqlBFcta7aXlaNqY2bDacbjqaye2rb8A4mF/Le/R9VYMq4401gs
06E0wi9YSSZCqeBNhe0yGvp107lfL6g158ZyEnlisZj7ThgHrCe27FmbF9vv44lIFkZSfTgiBOja
XZ9nOG25EMauYk+8WgmsSmTXJY/+Y71GFyaHOvZAr6hO8hQbErPGlTCBp0MQmbCmS9MtPXcA6r1H
GUKswmMGaYJoZbnF3PiUNzHHCEIhfLDKaK4vK2+M/YJPBMa5/x4fclU3Hxv4A6586uKfBM9XDM+g
n2Nyn2lfn7EHcBYqtdnheFePDgrjXTaL9J16x5qHe/BXJhgi3z/8vc5iVlUp08XAwHUmgnZoNhYP
ebd98JHx2XHRfZXmzOueM9t/8BGOwQU88Lja01GCJyiILXeKcv8yYxScD6EtxZ2YVN5IpNHmE0nP
woardq944zZJqaks8sWNI5JLFjHmTMP8J20ljt0ur52pHt1HuUhtmtMvb9hejopVaKToddbwCrG8
+4atKGhOSM2JWCgpL8KWSbkfi8yogtMyqKgLGElteV4Jo+N6vIERBLVQU33II0Dp2B8DBFypC0iQ
/XAW/qbqYfQmzv0Xb3AekaSXbC70vtVh997GppqT3KKfswAgQZOFk3ozRuzcjEXvWV2WpOd3oFmo
VBHhVPDi4HOl6KxyRW18k8YvEIg5YOP9A9Xcpxxu/yTSKeXmYqcd3WZA0ByvD7NVqH3xStSbjZXo
sWkgnkChf6vfcwlh9BpDv2cE797/f9LCMW6xQHfjhoUtvG+oGnyoGQBTOi9T29w/CSVf6JzF8IvZ
Vfko/u9PAEWuQqzRVI+8sqDLbAD4efaaNA1TeRcY0gdqCJinj8euOtU+ZwEE5vm70qMfpj5fX7E0
tPt7HHk3YkcnS4IZ5AJyOTWliuP/ii2SEQz3irdjnfXogOWfI3Bt62rEBK7Vu4+2TSDblFyfnRpB
x93axTx7ilmKIvOHt9f6SS47UMhXoD/hn2Ye+o2u7/kxgjAH2cmZhcJbMYSURxJb0n6uxVGAZ3u4
mkEuCKwXfD/48GTM8aT3zIpm+wOTW1/lKj3eZh+Qia2LfPPjZ1SkRzCLe4OiWaxe9FwP0X3lRN/C
Dsl6lUqGFBBm9Ul4z3RA/ZtSWFuvNpoIgwwDjBTsUiCfGCFuJwlYnvGHJwgZQfqiLcd7J41+n/j/
xVPBt2ge44ThUjGyNOcv62kOCR0eVbUbFtIJzQUs8NUZPKocNgqkY/DjAYJ5YRG4eFait9KUFqTY
7eKYtSnNVIhX/5vV5eic52yoLryh5Mp35iKfHOU/8cA1GhK9HkSl1PGOtYS5JU0pd8utjkOszKQW
4rBVPRdRUquhgWdB3L87RdocZ5FaXPo+SOz5l7BAWGJ4zqqeooTiL9us8BUU4VgK2NqBXEu00e0T
/3Z6R8293tJnhChaINd/IFNFO4SbT0e3RwbdPmxeVjLl4RwsD4o2vmpx9VbdgOha/FmCo0BMIDF4
jsoz1/2nOaIFxWJWJrJuVs6YZIe8zDIgHlDc4YX6SKIUFAOQmWbI7BP6uatiA/gO1oqB9BHMTNOr
DFpXXqBxyDVNVYtnjAp3czoMEZCkyPARUl3vuj9X0xMcdlRoI7oV5/KvczhXUcbsdkbfDbpEc5b2
wg8ahpVakFvIaySUL3f36NMaAZLiX2vqNNxgDmG7XazrnC+7IC9WY1Ncnhps/TK27tKpgNWmZt50
QlXsQK2CZfD3zH+qp05ak7UnvjP9T2KMSKooxExBJb2XmtX97GCalq2CbfQjAv82FuppZ2Xqqwfw
9SKfYMOfPQxSTUo29kdW/EMpfmGWA3hIZnzp6FSx+46cO97yafO8TH9bDfAsGeRREFkJruoEXq9c
Kmng715Pw5mIGK2YCihQwsH0mUeOFbrFbED06xYb2o8TcahcbKbgX7h1TyZhff3s/OB9l6l58/VP
nKwR9l2S4hqwuGG0L/ceFoABGEfIyBLP+dNGmnPskAO+q5xPuVnUeREkSnApfS5QebPiiKMNUB4h
Mb5X3GtLRGBT5/uCFCnR1FhIteYwZEZ12xdNoP10mvT1kzjSq2eJLD+5gn/Odl1CRjM2PgkAT0ck
r9/cq05bzPXZqDL3Th273JA0Boy3v2rE6JJvKeEpRgkKsZFfNSs4PR6BAuj97qtcRiGTxj6lDoMP
WmMa0FEDD/sRWV5XQQbqtQz43z7G486S6dbhckJizkySGSKYTL2ani0im8O1BUufGmf7M242Ij1u
BR9YhrEWPo9nlXO8Ckhq2YVSwzVGZcafM9srYevEBqda/5j3o4QM4bAZDF7I6i39BbEEdQlaSAA5
s5lH8lNl9tTqJhp2W/ubo+vOh2SfFBpHFhrasS6xZ04eD2xG/YJ7aEbSMxslxnOf5wtQQmHdaNYr
G6NuL7rV7N1TjnHwW3zNuT2v56K7fDIVAxS9bVIxYaKcTaCsnQhjbmkzNak+ndnERbrY6GQ/F194
94H3jo4UbfRhRSuBfbTb5SL93VbBQL217Qxx4ksd2Tymnfcr7cFKPYQQOoLBImhp578SCfR+Xfiu
JSlHmGjy63P2yRYVWEn0zerHfDazO995S8PTXa5IuQAw9mkslo2uuxGiHHDFG1YtcHjbX4geyY9+
tt8nozIF/W1MGotLg27cJ2R7/hnxQBWBemFGTxj921wp0JyOBZzcIA2q160hjdS0lDGWiPB9hX7p
EKPCPzUielhJ/oKS29Svaz45VRjLGBMkb5x4BlrKd0tm76ybmUeaFoL4zAGELnNZYRy3ifEGwfHb
M9ujbqe6iRpKGnE63yVcdOuTgG1AxWEstiBpjCPS7maDVtpdv2xQClQ2v+sPcHvqLZaJlTeGNnVI
Lakg34/03qs7CZQ6wlTk+UY6p+23UIxQbU1gC0M8PzQnW87Io8zuCZXo0LOfi3sYFlNyUPO1r2j4
9Osmzs/+30l/CONg32+TjbhJGPKnxID0O5b/Q6EDJ4aZwzwQJhCvrKRwi+zknHF3OXhMrHNe1Cn/
WjlJIMJPBc8UO/qg2gMKi3rbU2uCivRm9qq1ZitMxAvCESLv9n28UfvphSgXeNW9TgXHFNtywb9n
8jIXRN2yQvyH+7nti7mNcVn6IuXs7nI4RLI2ZkueeZJhpGbYXqJpRz/47xFNrB6y/Bx9KtvDuctd
kZr99M3CrfHkMI7Vvp4dqYHUSTZmX7Zf4iLLoTWBOJHaDK6MPoVl2RNnP4h6bsjkYOoiMWb5Sv/p
0ZPlEo15wIyOLDqPB2e9L3Frm7BBIUYP9AfJWQHHIZ1lNy52QDcIMJiaeXWpi902UcHUU30pfEn8
UdfrsfAFUAeAzL+X9ha5kDtWXpiTCKWycF9XW8uSPTsR2U9pI8SHqbC3nR/G1QaFzHqRCEGZAzvj
LfSpQv0n8h15qW2pNEEx1vfflm9yr3wDBN1kOTwnZwf3qnV3YUNbTMcvoGkB8II7io2rrdcm28zU
GeE1uEgU2OK/nJCYIFRZ4pXbrnpDsYVkp0mfZoKFwntAIYI+2/NVp4DWQxX+ZyBuO3HznJORbIeQ
WToQYzuZFTwgwvCLEGfKFGjmxeg/1LRv2QkIxVueQmxzxmE4n7/OaMDQNRBH5bpZCYbYkiMNhZPE
Gb093+PClLQGCawcjXbcgbTLQ4QHB+nglFr/CNA8grh4AsFqxgCkPmpF5U2ZjpdZc/VucGRiFl7d
Imh1f4qHPbTFbnSclSAI9FOHtu+9dm4YpxNK02dG3Zl3qlBr9KGhHMPE5UnUdBObr7TNVZD7QUMa
w1gxGqaA+VdV/gv3CulgFCNOn/86CPGx2pZvLfXZs5v4MgASx5JpBSeN2vc0IEUZuR9paZuGA9Ph
LFrG375YQhENiD7fbR37lluJkUDq2qHaScyxA+QRmAZhe4J9MEF8uo6ov7mfoYmMI3Ar31bFrTA2
Gg3HxxLrSesRn5ZcIAuS8/gSNvzx6jZ3NRv4lgtRh3Sd7vUe7IpvYQtGfznjqX7vZSO60uDAO78t
QsPbpMm2QARnK444iPi30AB4bIe7otOBuJuT45iCT4IcFfxkd3iK3m8Bkf9ErNdJQMA2KjqhSLTO
ZwixLDIoAFV+LdB9M2dWerVqB9Xth+rVH+SwAeQ+If0K+8v4gmSY4Gr581Z5W6h5FUdApO/tNxdN
/g9mnMHkXN893N6IMYsyjXAiZrFxs5ukJ1y/Ae/C4v1gXBXo3XRL9S/6xS6+z25iI45WDcmP4IK1
Pvsb2iz7vhDQ+mvBHwTE5wTVEQeAZGwr1jXteEu7spb3KFiNw7UBaFGali0k2476yV1ot0iq24PY
mJte/wT6ED8M5uJ6Hkv0uW9DZjg8bgXKexnDazi9o/tY5t92jbk6/nxJCMEdquzvCIkQn2isxy3p
GBJKOJR+L4+67heAq5BxrdHCvrxmPYLikvyRRtlulZhCePWbvR95gz2rhih7gWidbcUXKtyAwI5J
Gi/d4QQjG95ZpNFoZGxBD039Wc/lfl+huA6H0j08z6F9O+Ehlubl3MxEEu5hzloVKZ0NHY16Cw/C
MNmxHGzjTs8kxLo0TysNEd77qY/xY1ApVkpx29f2gARWBhasjGVigrWyqy7smq//x+IVbFvotKEj
NGK23r1zrGAn9Cxz6q8QXAypaQWA29OCPQMMc7DJh5kyubhncnEhOf3bZ/vIBjSTEjBkyigwrAzw
woH0tMOsBkGec+VDG+if+RXbnjT00Dh+jD1ZdQvsPp3LqQeuHXNeoHz0xOKvLNwfc0ffuSnz7Iz1
4mglmi+GX/TSKRJagG9R92w/XKvEXJcIrnVQbLzaO+VMfvmDjS4rJJ7lkf54MORVv46NU4S/jL/T
otqkfUVqtJTjZgwCu+ONXV0X/TfqjrjjItXXhNIvziAZGrEYkUafbVGOsdkUcgfZ8YutQvJm8hZW
ZYlkW3p8LWu+iNPoF1GqSFX/Z6cqa2abqE7MU2bAimps+W9BzLwH2nPggqD5nikULf5Up7eaRIT6
eIBemHi/u9NeyNFlT77gZiWuLwg6nU2acJEztQZNZNWoPbuYq3cJ1pMR2b6WIbtgpd+e5RDDS7y9
QApya1N87418e5KZJKHE0sc3lYGb5BE8f7CLFszNqDUaGfK9L+ZHLdFgXeihNvg+1dDuuNWFnefw
Q6CCp591W8Dx7cRuOlUjr+O2lB6TBA5Jn/zhSmH28Dh+/36/NR0O6rqdb+z87NqVMdkeZTUpsHQ8
tH6DV6wS+jTvA2ZCQ5znzpG4mP+VbCwaffr5+YMXkEEQrSUO0/KlgEb3Cx/AOr/qLOudeLvvwwxh
fAgIfsuikjavedotmjHG98vhpGwjcK53DK8+T1Ea07qHE5ZnqRJ0vdg0IsEe1G8LkV6vJbjf5XoP
yPjGFYqihjkmdtfDB4ZzRSk/sa+EAtagsC0bAFa28uLE/YlsFv51GlVvd2NekhJXk66OBCr+Pkfz
0FlxLNX4cWNX/iCA+EKW+izNs89QHnAz/ZcuymLZ6HEevkWWxfjaWAN68qh+1ggbffe/mhlC3mBm
OAw7gt0aSUOUT0QDVudL0zKb0KlE79HCMsbIKQ3P/L0sk4yfrDr4IBHh3MirEH81D7lWCVftFB0M
3MK+A9HhXY2lJaOCy3qBuHJJyHl2KDy7w5CHM+koVIz7lrKFR9URR0qAztNbYFISFROUsPNRxZuM
1jTqOlkWXJYLgeU1uPfJdKPBnD4js+2lC6iuVPASSBShBB7GqhhOeOgG6N5EYE7bd/OTpT3meIVp
MmKh1HnnZbQFjzbS5eE687N4Lq1J4xo4zGyiw2p87u+ljSYKbjbW+mfON6GeMSHHyEG95RebFU8C
HmNINS8V2fXP+IYhdWelXGxbpwwhn5SoiTs4Vtk1g00nWwghiSmNQ7xmAPKPuamjeTmYokTf70Cu
PKEPQ+JVLugQ7bmDS6ItcEh99pf+ScoRJcS61PP+yuS4fWwWHZz42SqgFf0h1BSsc4hL65Y7aGkg
QE1aakttLw3PAiTPWXFX/ikvUL0PWCDFUF5aXPVFRXx/SAsxGSrDzsUSz518LPOK4hmbcirdoNeL
rqEGy3jDFlVQkIqY6e+bD5oAGWO5cco0WeWNEGBdgEsfBQ+u+xLeMJIGfAxChD5pLNjSs0c4m/2U
50Nbs5i2wDh3NCR/VBPsbAg9zguMFLnWtsgNMLFM6ua6Sl/w7uPtMOesL5Ct7OcYmNbL0xmWoF9O
xcx/2/7JWq3hgpzUAvGqrkQfj7YJ/MGsra1DpH0OOxC6lgPrcZZhuWr4QwGeRGLB5KBzO4Vptm2M
6ig4hleAtu0Bj9t5YeFfmnKMn6gxyF5B6UTfUbVi6COADfM5syBvBQsdXaVHw8rCJbPONtFO5ogM
ebDdQ2YBlCeqNeu7+6CFpvhY4pfEw4wJRCMKnh4QhbM7vDDEyDZsMM9xgoJtcqwLYQ97HmnZLQT0
eevWpkZ5gJ7Wc7shDKAungij6bEBL/1+iwKll4B1L727MrmIL9FW5qMCw/1Rx00GM4KqKC4nJuIK
SS3HDIKM1Ha4WviI/NOPWlVodYK+BI3TIjnGRRDmCVuwy9VCEtjWOkpy6A/prLfNI0JkDXEG/OdP
eTktMc1+x9YRcOzH5av5DcGa0bAyb9DTGWjVi5ExA018UXSi0DlcB0SRjYmUg4dlOaRXCSX3mnkr
6GjoXLZR5Zie5DyFKg454V0PZj5noi1lHIPuF0ZsuNn1PfYncEhR6/g4jvBy5x8+0Bgg/xHHq7Lu
LsMl+u4dRB8lL2/f+/pQap0RZSE0kmD/dIovbHfjVDj7jonSpgNx2c9wIjDBn9qpCOiftsfMcgGn
ATgCCsCoyyrsGkegS/0Rv9pyjtGq6pUPMzk6Pct5wOpcGR0EZUN5+kG8Oc+iU4bPgd3MAqm1VxDQ
ozhwV7/X6hYIxC4wes2OEXLSzbKP7ce9XS+4/n0KiTv18pC5QPBF3Qg1vt3pscFYJIhkPaKGT/5W
vayu3i8IcvNTYXHj0ap8NiDSSoi60BjWQL26VJHByMMvxl3eZ63WkE6rSMAIF4MgliMQbEjJtQXl
bH7cX9wPT/OQYNU8x/al7i0BCi/Xj1ikHyXTquE8cb+it/PhXY8zhMpCO1rx8ujaH7yjaoduWxPk
/010rjinB2e0Q91VpJ8wCCCkPVjw9GIYZnp9+EKb7+dBKPa4i8VWfFfSif0g+2t0LWmOadIi79aO
n66P3J0nwTi9462NudCbnF/ajt3QaPJvf/pj4eoUB0iFS5l7BNh7a4bGsjGu4d50ks4n3hHt8P2T
WQRbtRIjdlG6KxPo9Ogg8v7QNnK+NQmPmokSTMBywg//8fVZYZCohNU8kMf0oDD9psDLawb7rvgp
bfMdy6+/ab7bZS7XTl1tnC8WnGA/ImuaCHPgm+api7Q+X/vz9osxkPOth/W+BJ3SqLvRPEic9e1T
Ly7IiS8/lRyp7f/Pu/D/EU2v1extVHvJkGA7u1ZAKmThwB7o5/AjVFYDTzk7x3p+YjIuFDSImbQu
8WPQUOBlV1HI0f5x3qc32BbA3rsZU6MqhHDY0XpJfxntw5+amlX5UoQMRHeBBcY+vZSXQSUsLX8W
O85mu27/YAdjCVf7kJqnibqeArBJ0MzJt6HLehvU03XgcT2Ji4IgDK3J3+TNZzn7UrWE9tva6diE
IgYecz4MLPFmfl1xz5dkGNHnyMspBaRPOWp3sawoQ4dYnWzzRrD7Oe2etXKX4u89IMCuMytID0y9
CziOhRreduUVxgClb5FAS/9X/ERjNacQUndzxSNwADfD329Mpssihhrc0EOzPudlLxwLeTfyvV6X
wmWqe7LoO2ypgFmOjwZYxY+Fv/Mljf+Y00IfbZq4RIOIel48Fytw9jVB3rH9PUDUNd0m6XrdM0pb
qfR+0Y+jjRsMZYSCDMLlNfrjHOZOd1+TKSx6Hj6oXhSY6zGAAjVZWJL04FV1DbIGN5PszgMBRDJE
Ey7ymXUzyBhrZWWT1rJYoO3/F2ak5UTJBKqS+KAnxQEjQHcfrWJ6uw/aSQmx2+ggwM/P6Rbav1x1
pQ4uQMhRfB0Ja/oFJRWt78JY/L7kvK1dzpRbjqtR+Rce0eW6eBqGDf86/lxcqD1wvwoO83U3PVBf
yOacBBIdl+w8zLKuZNcZpPfRMbPP7s6Bz0/9jC51hAlVcEG/AKY3XUFgfr9undjUhbQdSaexgf+G
Bg0YIVWmiuT8EC9tVMJWDfYodRLxxr52/oYjbj/RAV2OztYdDKOBKL7NewW+O85/KzpSB0pU/1n/
44jxjsf/zX9qTbyVJhtYa8m/nikFOo9eM+oAqrdj4EQlvU1Dvn7dOihsQ/qDhI6Nelat+YXtPfXl
lmLnu19OfxMg+N6pbntQwmuH0vL0qvFOh7VQxQBwsPYVzSCQ/tOZaF+ZEmrueojoThW9eNNUJuR6
0tw7qlRCRi/Gm5luL0Ni54CvU6u/r9oOAg8NPETiTGQpkuBHGIugfA8LSa+qpfEyJFUzJzoW0Xkc
impLDQCu1XBewwlVwNe1XdcSiUEYm1MZeB3lPS7Qg9hXjKueKQN2u/OzfEd9cU2v3Txzm3ygfoy7
eXQUwahmY+Y+TmZ9aJ89Bq3CMvH1uiI5YUnBBIc2GwVtIyDrcp8rXEQTMn2mzkqlN4Ezv+e00fvv
Ozu/cTkkjhdOKmFECVRmPYeP1yq+W5KQt8lnHNseBa1a1O+vbDJ0wIpXCwMe3qEUPp6CV568Ue4W
EpU699lII3xBR2UGfztik+hbEX8JeKUOOyF4vKCJssAv4I8kXyP5rtXJP3V97MI0J6GNpUFEi4Pn
dpZ4BsOvXllDeDwk9WebLOxHsP+Gms8a5fbEIHN+H/rRO1N49GUbe5H424xT6xbS9CK3bIQSZMat
jSuQmaCfMEIoKpSBgnS8y0S2T91htsSVGL2a0Q+iwK7Bnf8qrcIg2Qmw5zBC0vGJ7LTvpn7FZGb5
5HQqwBRBk8GCER0Hedf5DYWyhSDFrwjuycO1q8MOGGKARGwrjy4XdBlaNzhNCQeprx4tU9K/Arnz
A2flBN+MK5zLJV4w1Djm7/U6dZSokmcfA9gdNx1aOUO9j7rNzVZRJEGGGuxHq6/y7KJmBplV/rGy
fOtOJdG5s+1zA31FJHXipgaNiyOg2EP8/PiE4kji7uPdQBCRT3hpJFn9R8cUgAXR9Hlh7gK7kcKD
0UXUI3wNkpsVdDNzuH4/kNFQCJRQnBzn6+OH6Q0chMpViAaDevwWBPHZAejENb3tx8ypOGrpnyQU
O9+WO9alJbBsIotniEAhrCEb3K6Fpcokq/zPL3W0BIiR42sU67PJxknK9vKAOoTCgHYBB0lQL9u2
k/Pt079vxBRvoYfl4aZasblASiwYjGxzOwERKuwTjVNrvGrebFnzZR3T7cAk3MCH62mgAA0CKlSX
xm2o0HjCbxMU/ydZEiztUgT6RuLDEm7NpB0a42qJNV9BHdjRlVSMT9Ai3JqAUIfBj5iVaTNxGQ6A
8+sxAq9gyiXvJOPNnhInRz0vBFd6K0j7A3M62nau2SmndRsb3DH0jlaancQDpOSdjMMITSIPiM/f
ATp8TmvRzVFKquW7Pn9X+T451oUI23Cn8EFVmYu0tMgSdU3B2hqk4vGKNDk3gOVyapFtcW8/MrX5
kDkTnlzc6m8a1S7/ELP66MJUE8AuUM+MbphbMkoyK8Ym1ks22zLThQW9BYI0lv9Q/8GNs7eVwBPY
VPBC8+wEgyPRxG/XMdOmgYfwoZz8oDMa8fawUSA0GAUM5RyxP0fgRM0+Xj/YPIeuyBYOxyOI5v/3
e9gZ1lBbpthQjPkn/L//lspxfZkG5+XKnv4/Y1Bwcl5C5UgugWs+FIzBYLG6I/bt46DSte3XBunJ
1SOc9+lIY0kkptxPx2BfS/+mVzUJcyMYnq/LRp3TZZ80r9LjC5//om6IF8bRRGbdN1ULHFw4bGtO
yvI9kgqRGD8jzmuVnh7yWgNEz++Da+/rF+xX6P9ay5toemoji6KVXbiTcLJxjSSlXGKoeztOQcKV
LUbk4geD+G5ZgRDWVcw31QsYfyAXc6A76PbvWcEjk+j465m9yF/Sa+L3oGFcvCJzt86mJltZ2p5z
+w+5XCZSJztzYdiwYmR3VUdX3YJXISlf5uZwiFFsiyhSNYiz6RmClY928xrNEnLQBWzNM4DMUjZC
75GjvRilpSCtrqvoJCvt+fr69ewcLPjSom+ffceuvEVRt+Kx6tg53pSb7UI1e/SFrSvu/o/P5TCc
cs4NRAY1KllRu3muqrQSwTpOBlNuviHLN0sBO/X1dWKb+Bi7K7gSmPbYs5KKySukf4VhI+lFbY/u
BKi+dNgSnUzCmMmJMxG3dgeBUxPFWHSMmeb+pMu8/gPxHjDg8RreUwhdwgFgPIiR9oMEWdtsoSaJ
sjFHc26HYPTEJQ3Riv+Iko38J3zDrdoin2OvZ8IFpqC4+S0dd3h/aO7Y8jfokBIVYDIrUTytsL0A
FiSvt6qF2FpT9g6lVFAcU0Cj/4gYLCbkYJsrckcS9Y75ip1ye7kIqfZb862MNSY427Hs9wn7OQX8
+K0F3zGPxeokvNMolIf+fHGEl9H/IaatIm8tIx9eojHESHYjLYzO5lI2PTm6FuRkxZ3mFdhgyitU
uEN81C2C7hMN2pxBSXflEuZvW7GwR+rz51CQct4WZT6IqvO4MParFbkwpldMubV+hZdkDMW22bwF
GAvuUor5UXJR8t2UKlfCxBmi4lBul9xaaY7Lkkr2v1QgRCPdvMtCkV5uz65hBiPSiYftejuW5b36
wtNl4LwCg0BRR/KJmUUItxGUnOp455KEHcaHWycmVCOb1swIEVFhb8n57gDQyBOxm+TYg7TPAgS3
TXwJ2Lm9XBL8HkQWaYXCK64nyvyq6W8Q70ZNyWgdQBXfIXq3uzGV5nPeZ2oFD+skyVUbBwc9ZnX4
GmqOjfldiW6KbiLJypTrxKvOkEyA8uyKpGLMhqGa20a4X2rSFfuBpN4PVAmQ5V6achFbASVdDmQP
vXM+UfmbXFe4iDZNsQxzKDwmRmCyYLYTMM2J1hIBbob0M791u4NYe0aDAbf+evxTdDOpWT7J8QXR
Ykq0uuWbzVJpo0Sg3mqIfYl2iTVKGHEf6XBK3Qe6xlqBXVK+AEEzTlpsWRysPadBZdIeIvlAOR1o
8oinJ26KEUgVlZtYgFh3dxwc8Ig5XErR9Xfy2ENODpRTYnGujXlM61qysZXcwmJcgGZrH2ba14wO
qqYHgpfOlLCmwf7/VXLScgPNr9mJPRjOguApy03WciHLyUSPT4wMVrHWjwNr6rJC+qtiSrXVYHqL
qchyk72lX+2LN4nftYvl9xKHXnmTrQAioqadJc2kq3PEhvMhquqDPHlFaEVoniQv9uwpx0JTvSCu
+XxjOR+mlLixRCPHuRI2aEIXajQWr9wVxNLRuBXv5uTY03dju0cgqKp2DPBj4HXxI4Fi3VafUpxF
5Mjda6sQ3WfIS6Nm6KeRzQjv1kzETjz6qWBHU6ivdf5NEG4psZPX0wpopuxQL/fXMGeYw42pltRl
tqS21nTXK7uPLI1Uz47KL0oO+IvqTTfzE89P6cIy8effLg/KSIhEDw7h8Bd4vIKfI7C+GFPOzpMk
XghYjXaueofMQsO1QVN1rxEtCh3s+G0Gb8RcHSv/b8/DBsmLGYQx/sc8EQJNgNDiAgUiWN7zTU5A
aWIukHBLDbiyDb4EYjsTU6GrdGovxlp/j1qJYfKXRN56/SFU1SctejyQafE6IRSOei8P++dSdixr
MQahqQ5PuJEUdGLbW0sS3biaIRTPv3wAtwt01BoIcJkYFKcebIn35sZLcQGjLFp2yYwuG63fpBif
vaLvLi9VkgavBIE/n5WkwdYG1zDhp27wTzXWDl10I80WCqjNq5UZs3YtUq0EYKNbRe8+2iBSqH4J
rvoEtj72G3bW0B2YAI1rtSfSdQX/NxDsciARH9i/SN4Yzbsf62V+yzlE0CjeQsVdYGz/nBGUJDM3
at/pjBTW3RQlSI/mi3yaGoOaqxpDxza9e0truLpMcCVhi3TDb+s3sLU0BlW9KkRx5OI9GMDxw4AL
0LM++b5jgOoczDD9iA3uEZXEJUrK1h/PWLFMJW9smRioddY7ay56hkgxGW9kBhIlSH21RuEdHO2l
Nw1DmIsEXstwsnQx1Sg9zt6l/X0YPSK2ypmaXDtMeMYe7TgxOEytQAlWu+iXKFHZcTmfd3xICwMR
ldqjO1LGvpea3IHZBIrUyttMuqyW7xyHBv6KG3ZZL8bNOTeXzOC9d4jjLs/DIV/iiKXn9xW8kA3d
KbEFXpaiUAxd0oWwccxbJ1q+qo4mFf5+pgVdzua0dYXWtur2vUe+KvueDUmqZx6u4VCDvkErEy9U
h6wDNUnhaoj+ui3aZGDOqK1LSE6nq+YvozAAXRJ1qFhS33Ql7J0lQnFJ4AOuIqSmy6du0JgY1G/L
6EzcN42F72nbtZSzpf9UTL17qu3LiU3t5HEThvZCrjfO0LFRrplkloNshgrncMvx+Bh46bjNoNvo
oB2l/baSR92avtI3+EwrHT1YCGxK0XeNHXGgba+gc+uWu8Mo2s3yc7jgNojeaVUAP3zOTs0S3LHY
aQG0iJZE7x1W0WrtSu1dXVnUOT/jemlWf3CT0FKzgGtNZAdelhCx2YNPVoHq42HQFcd5yjKMg/rh
k3PtJ5k9A5n+r+EAkzHC+O1oC1w9s56/1lfrtuwsqH+HmWvdBiZZ/8YTg2xvUWHu+YtCEG83lfLp
ujxBmA85mXJkUGF0jkyQWNhg4xX6eDtiHPwlrmeCMWYA+3l0xlrFr4Y+2ni9XPzB/pedeGxuIASv
s8SkE8idd0KcGoD4PqlbMCAkxn27JqP8fgewIcctcMrmHUstSpv0xfL5jGeDT24c4Lf5gyWLfZRb
OLQoZm8JIjqa456nZNK22sK6ARYShGxw9XexhFZqeP0pXqybst/jD/oGxwxzVFPipTKRaWNZHwhk
ZrSxmYiAPUJV5gXJu0p+ka5IxohsZY7muIXIre8GwQzjhMppjG7XEpW3heqxP0IHHIA0aMOYQcAF
fb1oqvCbxZgtd+v2UgbkPPzU6u/qIW06ud/7xJY2j+jbPJ3GDAMCXQqFJjlQ/k9J+RYuwCGHxeeG
ymzFWNDtP/BQ6vbVYCAEGQyxNQ/bD4mSdnv9SDya2oH3/965L4NZsHneZQChXgqlVZqbhdyNgZ66
UNWG3siDaVRcPRViNxNAJZJeXNVdWZBlZz6b7IKpKxUI+Wiq3JyaQtVxrdOT7r2Mi8yzk9h75Nuh
XwymE+GFTEdWtpxjjNT5eiMrBmsNBeU5/lfVmWuVI4A1UZBSLfag/fSTnOe0piHgclq6ONV8a5TW
LXcHgJWiAXLRc5ovT41zD2GVZHTdeHM908rm4OhUueMQvcmYpHHk6yynDB0dD7k7yukXaVxP5Kb8
O55NpcHEGNUzzNQcgZQ3Y2n/xzWBGLYSWz+RiBbvf3HHi6rz6ZjE04xxZ2++OTWelF+j1UcY7oHx
UcUpXbu9Y47Z5+KTzq9z/2vzgitRHlo1ZPL1EDNKshReqxS8rpyQFchhZqcbuPgocCVKqgXcv2y4
25iI9hqoKYRI2peaRetK2eYeVRBmR27DgL6Z65/Ulf2DdVg27eLlfR81eBQflBdDF9rW1KB3WaR2
2+wGRcJxBAFYOKtpsQXjHwJ0aNHfit3QG3BRVWmCCWcxLiBsea5OtX/bx8gKSLBOIxQoXwh/PdSt
y3xQuTZasQFu7qatOkdVLXSCLtUm3Tjm+oP7Ou5IX5o/vfohUra9+RD0l0T26/zPABmL6FKReiNx
8PgmfsIzNqtUpVB5Cep+8JbkZe8CxYu5ippYCi4hDynSt5Gb+Ums0IR9OCFu8WevRY0dELtooIGw
W7s0PNoH6d3rsoIsIe5Ap5WHsKPKbUDVFWRjgAUlH8FvKGb48CvMuSXOjLnDSXOYgeCy9LZ1Oz7M
PLJvoJLlvbIXGkQZZZTr9Xz1bCSS1dMf/s26vafhkccQTCEXExJMbkSKT22dLavgvNCCuzlsDp2A
SMGtSIClybtEQPZGwVV/Uz001SQg4K6B0qltb63FhZpFEh+h9kECcaxitMrelj+NipBRCjTuy/cu
zfJsSlhbjvBii2iPCdfpIjqiSfl8Y3McTkUSFfD8KrG0jO2/lqZZY9Y0Ms2iCt+cXiaStMIkYapI
oPRWEN2XkOeiSsAppp+A8A+91W9xb1bSWqvyfF8WV8+UyZRmFOr3+2ZN4xr6cp9WlsdklplXyU+5
xoCO6cqBDFaN8WyGzZCb4GQ6zcQc6m62S0h26It5NtovMUfB4KGUKidiO9oFJVx1HzL6jhL/iSea
iKrZbk/YwHc+Hr5L/mgUc/TiZs71sz8lEc5wTZIwhg6y89hziL5rWnY3qgt3fU+swf1LryyDTSYk
2lk2LSxY3qqB7qafYpG2wN+JuT+k0r7OKKogX9EH4+kSGFyRUVtI2wJhHAZsTgvueDsNTFSyJ1Kh
egXbPoHQuWiD2YF86d31+6lQSMsP+uhFEnvcne53CL/hWjZyCPW/H9QWfg5dnYCVrlfd85s0iKha
s9AlGXkUwTAFl1xvuMDjarzkQGXTYfmFZvh5WrvihOWQVtqZ4WmEnXhfjyqjPU8lRV/jSJICAMAS
XpPzEt8HyBS+nIsLGCneka3cCYIAYpwmTWJcS+ENz9Te2vdkrqyTu0+Tc4J/rJbCc5NAuBDJHVhd
WY2X/soDhk1lkuVLVAvN9ENktMrw7TcHbLu5HQzgIB9To4QccG4LcnfGjUy/Up5IldIo+ln7xpvV
qdLMKm8Z6pdy0CmZWZzbv5BN0nZQZrsqrwgFxLU2XnhHjamvAoskSsccG9qIscNXMu0ZIrE3Z48z
hDYCtF2SH4JfRJafqzQ0QtamYnVIphz5wQdbl3ZWzBTrNiNwLJ0ZmUPZHUXauGDURz3HS+udNE9w
Z9VYwJyqSO6C5zGtsE2jC/F+YAu88cZu14VyxzAqIGkwlyPVr8VDhSTt9lDP5Y381poXevJSXva/
gJth13XNd7XTjcTSd+xMsTBQggxP1+DLlKhMBIFuiBOMmdNm5dWfEj3YTt914wqDl1syGF2B8eqZ
97EHmagXmY3YQp6vld4nrpErEDP2uYsfHeqETKI6Dc7nlJ56kqc4ckv6KE7oQUYjnYz0AM1WmE+X
1CMN3UUC0oowfbQtOjqbE54Bu5sMxcWi+vyBubLQpM8EJUxujdh9I0n7Oj1OA/EvdV7iT7BfmIeV
xG3JelvHkHzlPh7/xcqvEwGvjc6PdSwJ+EWJbBVRLa4LcNoALYqSeJK+E6HXs+r3i8MTIc1pd/xS
PJIO0xQqZp6scjUv88R9F3QgjTOB0wpP3qkjGZlYLMv2klzaM9cpjBpK3ZnH8uMf6v4IBtCk2E0i
V6biqO3zgtbjzQuS+dmbwKtf8GNY9Q5qoPN6Eo+XV8WzjIzkWqUbQYlXEwrQhBhabRsv0RNT0SfS
i/4HJCICsk/DejWXwF9e3Muun+ZF7w8i1Y44mfD9P1Va+D5vCrqrEyxb2NM1LmJVBK0Y8rBawhfw
kys17oghT3YGJLF0/NFRTbPasa2XBms+P21teBY3iM9wz0RixQJS+zeNE+5gVqT2EGWASPpRvrZX
qZDsJ8muLKns+R4IKWLX33fOJC8Igt5Iha934VYXdkYBlJHZCXKH4DPvjOpDiuv6sZ9XkOPM7Ixk
lNffBPJ3+RbmbqLIRKTiG8j7/dF/6/avWzut+3lROdR/AMcSM8mPFBzg+0LzTVAjm1hbldN12Bgl
Zty5scz4fpwHZj+T/NZK/Q+nLVE7glYjY3qIH7bO8YDFKW6gnG6uRSF1v7j/WdjVr4dhC3EzoVPh
x9feDtlivMuABTqZIL21REtsxICzxeRxXLV9LCNG/P1sFblPiIn0SQkiGn1PpVPlaWkayWO08oIt
0FaZlDj9natGenutIi/PQSNbDxKs5XYuuGqoXHjwsqmPKWCzKVbxz6wPXduS6qDxENBFHcyTEIKB
n+XtVLeOgbbp9xVSTZpSrgSFI4hrZX6VIEab5bDzG1y8ItsduLzOwdkdTAyJPdF3vojboyjCgmhc
OvRCGKp8cmkd+AGdugi0Xjse9UYd91TutDkun5fkX9mr2o6ObK5/Y0sl2gJC2i3fwliDZYWcNfMu
eHWCsUX8mAiWJcu5OY9gD8t+1SnP8/pd1K5y3PlnRQJ26hGdKP9Dm6d1cn+gyvhFEKHqY4N/U++9
0yra/UjaOGK2lpSPOUsDJ/qgKoLa5V5qUmChB3P1Krs8ZxObBTyYOhjZLkJxUAd9gyZBcYrY5+5c
XYHWoPFgOVyUazwSNuB0gO07QLjI/yTvpuNnyo3lueLj0ojifipG+TUWg0hpXBXFNYn8MUVk+nj8
UNelwiOcgDGG9tK8t3AkTZQg9jjqEG4erdp0tHeArzip+OdP9/KXXaPw8r0cX/f2nALOp4UZ4rAH
nwfebs5b/soBSFhpU27myRzbl4pLgRDMSm37qVV/GceRpodPC0Ttd/sGkbgs/sNiCaoJJapc5biN
2jFtsP2Kd+IWElqiAl0mdGuu6ZnEVMGfyTrXVFge2mlJZuNx7+zKMKSi0PMbc/yMJ8OTMAUSFTVi
LdIfqIvEb38y7AVGIsw7e0Sx7iGgmrWQEQGw39iq+JLEhN1tUy++kFLmEoeS1fukeNSnrKcXvulP
8goSYAtuBs9ibcWmKci0UcLaOezztfV5/Jaw0QXFAV32fBc65+SkxQ8slBOqBbFJn88BH7qi4MbR
0eV3NGArXphxhu1w5aZ6uNvsjba2UWghZ5x3c7R0M2EeVxL8mRUTZvUbS/qZQnq+xiy8T+dciRna
CBkSiCnPCjqm+EEjHEfQizYn0Aw+LqK/EbPzF3ZULk1mMSKiysGPpVjZ10emnC+7EeeQrd9WyJKK
1sMjKd4y9pDyYvqpbvUF3Y+zn+NawM+hFg9F/+Lmf16HLGA0iu2Sny+X5WdRCjAu6USV8wcOo+Ee
gUSwc+vpRQzQMHqqerDYdBe8ECtIh/3tkqHI8asLCho0wb+61UYm1oszz5epsBekDFNbIFdwq0ik
omWTO1z6oo87+7Gz6Ky2+GjL/zBN/JZjXhPq0mBLH2ZeeCYETzrntLPIacVHl40+X+fZJ1b2k1o6
YonWmxpLcOisRB7bSgNzF2fcUzBYS2AcvE9NlQW1ACAELoLW1QwYIve0cgPwk1dd0PMaarFxIlyb
w6RAjZDXh6C95y4mY+FXd96Bg0dOQFMV4Vtuo1giD3SZJo4faWbw/DtW8iQ1ET+LCELzSDr1A2zq
7ATY2P1ORw1xVp3HObx7zhuxLwgr298G6ihpesLUYC23nNocWeOiA2YI1q8HJG9GrNJK1ZD55D4V
9b1fb6ZlTH1acYJ3b1RP+r23BprnCN60pNl7r/5pNeet7/nDp9/cf8hR+iQMgfbY+14ZcVk9WJry
7pcxc/ITflXfXvsbNclAuTSUV07qzOYmYWirCF2DR2oUj1J9UoaVQTD9CYHfuN9fCtPEb1mb0i7u
o8B5oOtWUPSvbOt/h4sxqy/0tgKz/7LolV/RwoMZ2eWRJL5q9E7F1p4IR7jc/LNwZwgBCPBh14R+
bZU6EEkRLXQK93fmXSfgXbJJ5uyZyfxYIzrVbuuRpr/9Fjo0fEoeH+AjGSdPSigBmCvczfk9Clkp
hBmWLplW5dUY9DGTSTqTebpeAMDvcSli9cB5tMndDC4w1OpphaBNgrumoIEq66zVNskVP10CfBCN
bCmWO5By9Q7yLU8Q6hH0VFHGJFPq1M3wai8CRY5qD92HhymYLzeIEG+LfI17JzZXkgBBy7awU407
sy9zN7Ll2mTvL0PnUo2X0XhT//HOaEXt00wh2fpYF6NLTs4wS17NYPLscUPyR/AsPz0208VXHxpg
/zxY1TN0IfCT4WmuVgvolPyOzan4X//di8nQ68NjeXMvXXItyLMzqB/qJgtK7oJtk/SiUnPcMJq2
w7y/XSv/09k9a4LSn+36N45GQlpRzSPGxcY3ohVd9LjU4bB8jQ46f5AXB7S/I++da7fV6XaYTTsY
2xE1iHLi0mreWbLBEdU2O2UVkE9AN6FmWitGFX4t5xLZaVGDYGoaytAhuLAYuC3pX9TZ4u2gZ8MF
9wiXpeLWV4RCBcULXM5ZIIWX8WxQ7E793l0/IJlb6YF9AaSn28FstJFM6YDD0uR729MJofyhVheW
E+w29Tj1U3/5qNPDhGIoS5ZaZe0TSwn+PDe55L0EIaq3GnsKX3TVzdgo72fm4W4eWPN+1xAQZPvY
7yrgoAxwvdSo624SbApuj96m0ctfe2kYfIRHd7lXQww4cJENR5NLoNwrESPI5TDO1czS5Mcrvl5I
jIv1WZK0Cu1e5ccvwFLu7WApPORmTOo8yaNlLvzfH14w9o4VfvLYpaUeSyVVyJYsZcfxi/2rHMKU
AtVIp2m++g1nP20Fl9s20+xK2ZKxxqBKP0Cqq+SN5H+sSxQDqfiMd+RRfg5M0yA+w3HMDp+HQNB1
g+pyssYVunyhYCn26hq8+TceCXRwY3NlcAXkQy4T57dDTaL1Oan6K0md9Tmyk4p13+/Ag5axBiCG
XcqpuVkeQbNAF8ni9OJ5JLMdC0rPdV7qLpSx1EsHJBUVnFCHSeH43pmNefi5OX5U7WWNoY/x4ju/
/qrKFCzcmWcfCwD381FXQ7r1wd9DF6wgut+i7uCLx6unR4YoGvb8+GumQD+/aZh9nGiZn5DuPnKD
kJnOg6E809V+EJgKz8003xutM2MzIz0EOZYnLpheFam0N1EMmwlS9Cpu75GVAqOtFS8Hu8aNe+0m
BD1tWzApmQQUf4keCYvX8nLrFpSFB9nnUlWYZd4j8dYbGh5MxxkbYsgpq5EHopy2UV6I4tuP6kCj
z8o9ggZRvdUKhhvFA3NYLbU9qeaIPymKotdR3nPdeWA5a217cCE1AS1ulD9sIvBTHs5AsS6/h53v
CwlYXl0AlhNZZ80C458VcxtrVp9wRS2XV77A05TbxpPWa0dpmPn5RlshsjTyhaQ47Uy0PtdsJGbT
YW8UeTyhKVpjt/UPKpJ5bs6dRhAkEHgH3zFmGOJrbCmpswEKr44aiz+xBwQ9quYM0PTsbPd+RGsM
i0WlXjyyDfaJd1+R1dzx/7fRXmF2bPJgRNQhqRhTFfwVJd4q4UJAfxIkgXyznZ9PMK+ytm7VrcFr
g9FjLOMsMzTpNpAlHTRnNUmjTx0bV7nAEsOvihdqU7bgo+YRxRAIeu3GKCAGuNjQ1x3I1JkrGDdx
JVoTWIpIOd48FLMR8dut8pV0ujNi1oCdM1C9+55bzgXiB2V/9AS7lkZbVHIM/3+G/HOQSIcXiaBo
qI0VWEkov5vqFH03pGvfx7WOIJ2kS3rs8lo3L+ydR+AEjwr48sqme/Huf0GXhW7+h4jbYOIjvVDa
6LzsamisUrXLkxxhu0kVTOTGtogNoGMP1zjY8oV9wlQWDbRNwZxit7rv7iNe8kqX7xc/I+TrwJY1
/yM6z1gN6XLn5XMVX7ZzJeohwoXq88dmURzueRzZaFQe7ZwWJvbXuCXv1GrMxGkb2bh/4bp0fItb
MtLxVO3zKx8X0GtQIe5fb9yFJBKDRvpI+Jz9qwlsbpES35oHCz01Hs+DWRbUm//0WJIHYPnMLLt4
TLYQ36vaJwV4hPJb5AWPZ5RejETxt+QwFNoR8qpWyVehgvwXP1MZqLT80Nh9Jb4joxMz08CzO07a
3xoAdglp52FKV/NYI9TXaNGlnIvKlUniVQyBH5jUow3vIwV1YugYGUsbGGvtUhPK5/sSiLOLU0XN
zwM6BYCoSsa2DFuA4fsx8HfEeDmz8T5/7gdea34LYnittbBmHHVZZ9FaicAkkdQlv7uWFKZK2nKt
dr3LsQN944KTtpV7ihAKM1Oax6H40f279K0kRSoFdjWmSWRWjyCsoG9mlhbgCY8QVMu/eb6DjG8Y
eavsHjjtH6E0pcceiB/RRTrF/UiBU3XmnPJujUoZFv/CmfEYF/umaaBx0Uz1675uCXGawBNWbdPf
b+ah5p8I0t8cxYmtcrDO6OhCmi4riLDjLf24W4r0fzau78OOvhLPGGjyvJH8y9XoS9d5dYenjoIA
9PrN15h3KYqT+7YLLa1TBflLu/Ts2n6hoKTwNJxC+MYGWv7m8eFDb7bJ9Ti2vd1UnGNSY/PZF+El
dDl3Bsesh+mK67ShQf/ynoqI5CcHXVdF7IJK63wPfDbmWh1GXlv8M8lkGEotDy/aP+Rn1fv66jQB
6vU3IRO2YakMTygD33iQBlWbXCRkuTYMP1TRYHHFFyXTYJ2xQ6PCilCH8ZusKNjLj9BxYVebb/GH
S3wDSaHsUDEYLsAC6vJQ/tTw/BbRBE99znrf6z3i31Tfg+EBrXD5/lJAWNC0HKRXj+H9h81Y4NTE
uwDFg5BlmtmO9BAFfn7w4qMSDZsXbjy6JyV6ehq/WDxiUt3goygIxmPhqyjd8ShFDFkNHdOKAHFb
Z8HPJAhlQX+U9GwReMO8vXKNAbgeIcMst8EEDpaA+C/vqsUK8wxkrHyBqvvYLutNxJaT8M+9TYEB
ZFVlpdgfl05wj2N/czzns5qhF0ArLdZTUdaFMZfCZnPePSli7ZLZD0EEb/VnnU09UYdjf3pRsaN/
ZZmDMmyHhVjnUDCKes/98EKrFlDBKO22ZISu5KPRT0KrecDm0NB2qlb/jQgvVCkLcghortkMY4i+
zjrmV33mS7afxYSdvIBBB6QEEDq6j37Ql3MACNZi4IsfkJHt3Y9EMP7Wc/9mplBqaXDrfAbRpAQc
oXLtTCB36ty/c2DZQuvX0VHLYyadpulnQ8Qij7/dRgLY2vv5BTq1Nj8OZaqRzPEe5n/TvR2OK13F
sVUBMHSR0VmTizUkAu6OwrfKVCDWySwMUJw4wfNAbXF0OZjChu/JeR61BfIaGupSBoESFlyPAc++
wGC+IoGQ+LSa1pqHxpda6CXKvAasJOjIMDeoS0FF5OZ7jPfeqmKJueRclp9sZaEuIXbGdP2ygWUz
arzUMPqpev6IbM6wKWcgAb0Y/YPw8SxdK+KSbgPClHPGGqZvYZxT4cB/z238Oz2xcBzy6cJ/28vJ
kSe9+RspIYPamrIZKjOtdKJti9cLwUgoJ4pB0Cu8PAm6iV4AecEczxiOFNb6C/zFHGV5FpdgZiC/
37rk5NgLjkcLH2yTA9VjUxLX7vLG1YcMYoN66gvAm8yvMJyHoqFT4Lzm6d7PYlkGSdFZm7sMxzNp
JMho5DJTPxjkxzw3q2yZ2eQ3gyDn/DrBYUAjNpCUMOzZvWVu1LyjqxOcZucC6UjvGH0qG4wudARB
+Fh4ttm3E1czuM1Bqx76okWCArLDUGipyi9x9BmCEvtK8s7uC+J3lEdlRwfCipxnIPKomqVkfqN9
MEYFN6yxM7IrOjSHRWVRXO4V960CnGubBhZ/4lfM21wGbV7jPgLqSuuYr+8GHtr1y06x4rX7gY3K
9dfMPy2cvz7i+ipqXK/N2m1HX1Ku/VgpsHmNZ6S/Ixsk50ZOHmF33dUNQT3HYdyMZgPv2gjxwHtr
Is6emZKTWxx3uo4ouOp3Sw6bSgJq7LVFMDuT2/ZMplAzEi+RDvDu/0G5pGSGm9Kxt+nUOSeGlSRU
0ub7L5pkJB/ywsI5DWpmpjVtRdo7xjU+tBKo2UYtM+QGBv+850OCqQfi8KsGIrPGUsWFuG9w6rZU
KK56Eo8ZVfkQD+1mvNOEjvl679A/oKNFcZUHzPCz2qdik9dU3b+CqU0lGCp1LX47+bu19gt6iXPO
OnLLkF5X/nUpUqVpG38yv7rYcIkeE+v9qZY9o8fQAOkrMwgJfB24AX5pbNyPLJHmKz+Bh3kxdeFo
BAhjG75ON+i66AU7oh780ZpXZgQCFAtqjx+zietv7NegkPQQDKNDkACZ9WzYIu93naPQq5Bp30tI
OL6XARpdSt86HS/I87Ty3miMeQAO/5TXwGKMtAAxRBRnvvxe4QpxMjHyxqaShhluV9WROzfzl8SA
IRIu2IqH4BnDhEgN+cdZY1LmVXv31B5R9V8XUun5lURmBda+LbvhsMtGOGZUJYax+zz6Tz2EFKMx
ogGg/u8mqyMRnNme7fhbOiXp+yqdz0VhZylCM7qbtEVXt0+L7gBkgHVsIt8RfJW0UyP5OyLQZEkG
dLNEE6a9eMczUkE4MN0f6eSareunrsxoP0VdeBrwyyw8dL4cIMchVgKGxA30Fr32DOkBey7cnjPV
VyTFgO+pjEsMX4bExaClqicaGo2OZlwr0JbQgG61a4HKYhMVOomhezQnA4Bss54qzTEJ18vObTHd
1a1ubXHs3UyB0eWKdwWZnB71fk0AlXTaH3eeVrEQJIdpgLChRMiY9KSg/sCcWeg9m5hQnERij8rn
oFWDp8RIklR4gPOqCCOzVkt9BIaxQoqk/ChrxM4uIkm76ZhTwBK9Z70PKH9LXjly9RDwS+gbVhML
twt8o9DtnQxEp+ywS+zwkEFl636q5OD3lr5v1EQimd/ge5159KokTDFwTyuj9GKfFkPmnmRp1P4m
Gl86It8bYvztUON2H5GEyZqDxFIki5zQBddBx5CDgcjwy2JpQ2hLeGHOMRA0q2lVEJf2xX0DkDHQ
IdmZuCT9mN5oSojiOpKHpG/QhfsHFjXlvRZYIN7humXdU7rNjKIaC0RSZUuB5b5yty+F1OcXwd4/
O73bzkbcetPy16ufkXx2weYiiv9+vs70MsEkc7vyCOap5dTzMnqhZ+qYh/x6wnsMdQLPxMTogOC+
i5onaekl2sr747uUBRuBp8BFlRmFaDh0E8VLoVUB0dvrEBmC+vr3NaniJlHogj80DJYSewEH+AJI
S2dEOwGQuLjVkk5zxkXbvkflC5nPiNeF2wPfCUPjqizBFpqpcDNZKjLHJK11K2q8WTc3pXRW+rhy
VmPq6TfGENOp6upRlZUFku3+iLtwMM+DzGQQQKMa8SOJDjBhS4rUnBlIoT7MgUY9tWvrPFiX7i8s
JIVlX1t7D7cDOxRWPnM4b4Y3ijplbdQP6Lfj8lqMOqJSEM0fhrtBAELIfbYA7P8TQsF+tBz6atzh
J9792IURDmCVPpSjcA4NWtLzUWgOGMoEAmCqkbjq39PqmbmIOvpngWjnI46gCVXZRyJtXeyVm2lX
qjrgFdAqhbXuucs7EF+tTpPEn6HmIrZtDsVJv6F6gWKpsLzTS5IsQUw9ZCyd0NoGhSKB/91W65Um
V06d5FtzOdHOJWq2IUMDuCFmRNMkYY3JFEWj9+3ovAc2vmv3x8d3OEoYt2npK3wvlD5tDOlOuANh
wCIgUDLwpjKZvszBuPRaXYxfuq7tY36bQrV/sqTpY9Wi1qz3DVfuumiyG4Ei3/GNAR0yRN6/AOY9
wfx9mAOyyBggJuOIoCtYS5tqjB57ew4rbK7DOmuTyzPAAtvZdZWkMRuPK8VFty7nv41jYbHbr8MT
Z/oMzE2wK9YAizEQ2W3LNRHKkWkRD6v+ddlWE2PN3PoTcbuGaV4SwhbYhoEaLUeL2Vl+tXVDEYL/
GqtXsbZaPSEmezo8C8QuDxDTiZBGdjipocDVij4R0QyGoP1l5YvjAZxHPOpkyADykI9uRIlv0H/h
q+n1L0axxPwHfqVakxg6I/Cv3hxv3u2scnYL0ww2Ejjj/vGcJ4jpwjCzfKqGv9jQ367pZLd5nTBF
wGr3wzzLtvfhnaNGA/NcYvOO2O3JLXT2W6B1FCgybJ6dWaM5nVxnt8seRjlY17yr88DyKm/tpVDt
L00bkIEepPADftv8rfSkkN413txtoJD6g7PD9LV45a29R7+0QAkC2XqF8yqgvotkLv2mNF9RJSEM
tgS5I1YSGPsn+aNCTSCl+IRGT2CHSh3dFzCjVLdBJwtudVv8KS0+NWOCqUC5vZLuPNTIo1jomUMK
GMbgVTTiFmJAs/o7TZxCqnBouP6P0MXmEm+XUXTcSchSXZ4K3YBEIExEk1bh1dLlbS7B2Iw+43RZ
uxUWwOvfkBE74P/echsSf5Ji1YO0Ad4UGyDAIP6B6RGUfnrDj1n/UcYkV5H3jgs50HcheeXz6gVi
2hA3lS8Xq6MIhkMHsEzdztsHmbESrt0/h2cPJG9F4Wmmxh6NhRQ+81tWv6LvjdSZ2vgnvAWl/yXv
Qq6ZoG8hE2w2DI/Y7Rw9oXCP+whnpA669ybxCuGszZukwXRn54/8DImiwUAPbAWuKV5W5gB5Hx5N
0HeR9BwdTIIExhzfZWs5TJkuoANx6vdBOanI1haEDYhDVvZmDNmnTp2vSqlYRv/xLVQPGVfr1yge
jvWjhQAmn/tP2EpJ/XTCE5J6sn+pcMyL25ZPpixcxZSTQNV0Zg0GXfoa0XbGtj4cAASo9Uu6Cnd4
Xesdubl7s5EjWU9eeSNAlpgERt3U6TDaeAM5wK47a2RFRDTl1j7hYFigr9nfL76X9cCacj3PCEkE
vaTq0vR4DfmESscZBTDNL871FA1dII8UMUFk1eLbjHvay6VqmF8VDBwDI09w5XyA6szWuN1xFke/
HIM1TTflS1pfpokt9kN4qQrN9obRhHy5zBfLN4gMAJZ/t73JQzGWIOX+mXQt16+WvciFDYenGBJm
ZAO4zTEqeJNpNlMjsGBV4bbhWEBCaLPRgpAk92HkhyR2QXeualAzWjm5oVuidyKilyDga/NteHVb
sAnBnMC6xe3I5sMSnKdmelKj1Tf0OU5kXQAtsGQBPznWE5d5jup6LIq6Asi55C+/w0YS8ExcytN+
7imiYwh+OgwYlkx3uycZ3Jh6c9wQWbg7i83Y2sSxGlDgT30mxAZz40+cISyzPoUxv0v6GB7kmRAk
wpTeH10WbD95N128HwRUjk2qzzffKt7Am3cjrthgHuseS8YIxEm07M7KPkv3BIr9lT57WAEYcx1B
Uijysa5hkVLPgZTcMnupiwULGQitr7b/zaQpvZXrxOfOlajA/sTyZUJQYXlY48sEU8M20Ni3+jRD
5j3nWF0LtmMb5AqiuEpqfdMHX1eg+P/zyO6mwBb8KCGQ+HqfALi/OFpt++WZ6edA8GTvduLIZrdg
y8pq69GpJ0cV+Bqmcs1F7/bS8attDivBsc2DTaCyXjiIbNtxgFuKGePsSVEbkg9//SrRxh/AW/pg
1ZgnIWN1qjtCkcclbdHyy8Z4x7Q/ThFH9+XRvTgw3OiMMAs+RzeVVnsXvrE9E11zamBC8PYVeB59
ZluzzCjNjKR4bioeFHUmzt0QM0fJkieDR0HJr6UAHBLWLcUkUjO3GWPlH3pvV0kyXOqJ773jB53t
/ZPPBUiz7pRNnA+6eMpA7biItOyb9+vaTUfpaimHIzs5Dvhqo+aQzF9XesNn6sCM0PwUic7MuIAC
YP1qRyLEydDZZTy2Mld9pOAsTO+hHrPApd8JFSNjfKWKmFyhqxFof4uNGSNvRMKci69BsHsem+Rw
vk2UlYIEaiFVILsBT5b8u7FuKp74lN6wn4sUIfG9X6wA0NvVv8m1jrTQWcv5UCLrLraHfTD508/6
Y8n6oYd5tD1SJGMdW8ZIkPMfrLOjiTjoDhGQG1iwuMC1m9VjkqQW07IgPzdlU63XaU4222/vlR45
WJw+rRDfPm83UK8lB8get1VDY2zSeJth23U/n4l15eQyqV4rIS65CT41Q/w4OB8/Gn3QSKVrG1n3
PUWeQc623ng8ppxACfjfRMgEAvTQCkb6ifAOS/n+vdCInHA5a5L792v56uS+AJKxai218gxb3Eeh
3Whrz3Z94lP4ekEon9dIql21cnAHzx+3YAFhzzAzHg+JIj9aFdYxB4fpXSLkfJs3K/Az90WOK+Md
u7PfOxPYDNveKVwCFln+8LavclC9tvgT77AEM9jjXEnybM9fqp16TkPdk9LykSIfD72k/YUHvQyI
okbimkxpDCNAwACGyLGFpNPNOPzV+poDQc4MGCNy8g8rtyun8SlGN8VZbr0geBXUtxMgcZdemPBb
kytWzleaZuF0WTx+mPGlVtlv0da8IYzjnujoAH9qCOIHorBYBh1D3wTTmJfkbtI7PwD+VHlZS8iI
QwfyLbUaWxfDVEamqoh8aodFYF/s1ZeflCD976xsw0pPs/5N1FxzQvDgp5F2w3e966rqSRM/jAOe
EosBUwguu+Xe0WmGrG3GaToCoG5oz/+hKHfSWmOic6SnSlTlDS7h8HrlFtfaEcwIubZoSkqX7xF0
uZwbYpwEVf65UoKlTGnw4lIPu5DHG4gV0De92xAY/0n06636r/wXKEnDEbDTLT6FGu++DQKFpUbf
5YI+4154D302PkDjR2jgbI7skR9e390N694bI/x2QOJCn7ajVL2ZABaUXUIrsvsCFv2mjOyrn9iv
C0mvEmcvxco+LgGTiY6wSP6NiVWDBfzx2kdN3rOIfa/LKJ8Biq92mLQTawx1VsKIfaNbkOi5AsTS
UTb7K2OjSL0ZLLh5QJqcdh6FshTCFp1BIPVfGFKP7nMX7Ac0dDZROCr7L9ULJdUX4GG/SNdwbLyC
HZugXJ2afZlXRjQvQ2GsgdHltvgIjPSQK91BYdRp8LszbOe6yCKf4fY+wWkChaIWjd3aOHakbueA
XE7Z7mfD99oZatwBVOnNI2/7lGoVeb48CLnk2G0Q/bQ4yYe666uWYSxHvkvlCo66em1CmvG/NtjP
V1WRsU7WoSML0i8cRlXUsK1wuqTA5p5/wC8WwW2NXXF4Aom6UexfdRcBemHCR9dF7Lzmg+RiJz2Z
dGtIXd9nrj1Og5Xt273fiiy3xNklgFtJb7HS8F9o5lnRIHx1LQGwlgZXJpKF2kKG7yFR9zW6TVbz
43EY1XmQig/3c0czyZB3+Repw3PYSJ91/+4/vJhPMUTx7kTrsyTwCidGYE5mFSXge7vLZ6cN5tfs
KG3XzCfm/cgvY2QiZ26B5C1vZ6oDo5UOROLRh4YIbUQ+crtVJ1JzJFEOc0HP8AuA7Q8pUYB6IvcV
MB8LKQ4cESHqESi/I2Z/HsyGY6DiRn1MaMiAw11hiiq6iF9l5KwW8/LwoN+SjAguphl4qh5M+zGP
rKpN8imPelsl8tjkdnsGbQBWToXT6hQ4nBUtRfMSSAuUrhebNQ4q0dJJQCrIysQmXx4GwSzPoQTA
jZLAZRxdWmaH6uLy9jofjinxamYJfb/H9KlWuCfDvkimE/c8UYDzimbNz5gOnNkHoWl1WcPDqtfq
fqA4cC5Ao1Xb7UNn5O5OvvsVB8WC/3Qr8inRRosywruUVwRYT9xzZ7JN1YawUVfKGIjvW6vl/2hv
T5O0r1KZMcPPd5K8WTtynohAfeqnXXOG6GF6X7231h3xnnYBBQeoiRRTVBeH56VpKCUttiD9t051
yjAL+D+oSdvIpy9QINPsYqrZThVt5LLFkgOWdguqdqYOUgkV4PHE8BldKNMzWHdeu6k6tEyTWxPy
v6u1v2wJxJ81IHr6FAmc9SxHyDXBbv7sAhvBDqQhPeTZ4fYEDfL5WrbL+2Y6IB3zkUeODTUMZCcZ
14LhZHnxfCd3rUgTnlYDQGL9fJL5bkAA2ayqFs4Sgi3BlIdLT6KvxU1GiBaGFcHbhJOwAVBAXsBG
+sIYAjvsz8Dwhxo5LkkCCJ9FuqpIH7g4oDKdqpE8YZF9OFxq+IrpG5Y08Qs9xGMpJzL//7FVGL2i
FXQzd9tA2JqBXEhU7wR+/7B/xbX/78sum4T5YBMXVcy7eTUJhC1Iy5FXiT6I1m72SJllymGs5ltR
XaO398Zf+QZahRJ+6xj7Chsp609HKU28HVPIPXKXd4+9iLp2Yk9+44KAMjZibHJ1PBNeGL82NNpl
EudYRtMRUPzsYeK+7N/HgkpsPspAx6vpkCaMsosiLnnel1lzwUzkFTQbkUVSG2eOIm2bB7vjNZ4c
pCR9TEdXQn/HWrmkeKRHQLTM7ziodWrkH+uk4xZLXi/iMInBo84oDeF0oIENJjxfyaNWZxCNxaR1
Ov2FNa+7p/xaKR3TiKSKJgjnTIDjl2+NnEMrRcqArSChy1Ebq4uaFo9CwJTOaqXiO/BZ3vdzHabd
Z4gPBJJpzvzn5EHMD2SrszRxxzvVBE7PW671HNKtgqjYpiYurO6zviR5KN//0OGJZfSS58BmxCOZ
6L+N0mb4WvD9gN3HEZPE7BvGew5QxNt/1glIa1K/Bq4qdR3aYzEGP2iWVDHbDEwUA2WlYJlk/BJY
mmnpkS/TWcTlyA7ZHzewzrl1RzYKfssBN2LfHN9MSZWarRBRHCav+wwt3ajKpVztqIego8GP/nAs
lHPI6O3SllUNadSTjFUphsCdGee+NRl9a2nYrt2JHFuMUC62j9+16S3Evsu3OqFrouc2Q4MZCczi
iiyjUwkz7EgeLnM6jRGa5/Kkw1A41zhvxLWImq+Q9RUO0QKRlnt8BnHwnJoN7TGQP3Dm02J5DvQj
n4hDJgAKXlHyjGaCR0KnJhGi9xl6Fzew6lEmlVBYB0B8Mt9o6pjfqfqP1S+iyt2F0z5X1xrd8dGy
IfikqvBqMhMJ+uFSX/Nvk/Z/HbWT/MhBzllfNDQqdf5s3qEGbMFR7sMRE5T4q9uNzyT+TgiwqMwy
804bvZBXx5qnpimu4udi5f6DyEC4pM1cKtN+pCHrrdI/Qy6OQg5UWBm19umC+WitaLTJtiKpcUbp
zXggz6rDdkdSL3kAEdfIK2wAKlk1uommZ5o2z9FNgR3llF5M7mj6qCI9L6p7wUY0BGZjIf3JiB/B
lftNM39/JrJWHojWXsKwxKqfRB6xNhs9a6hBNOFWJyA8I4niTbLAlxVyUP0VS+VveADUs8JWdON2
sVXtnuT0sQ5PlnuiieXzVNGIeHmaoVZRyv2GsO91Zm7uJNpw/B5qT1qXAVh8NJEal5Tl5F4ziwdM
Y3BU2TPDu1WpZciMOUoZnD0z9nk2jgJUIuiVvXKV47h1qtBYQsRbu+x1dXyHo3ujoIkBe1Dunah6
Ib/1wNZCTUkSYppSHg30tErYZGKsf/jxlSJPuyOd1gLuu69js0mdeTL5ghM03ciXfgdnt2MS4FrM
whmY8jD1rEpohLlmiOzInRRgiAlY7OHDWXDHRPg9a2nYijlpHn13JSZYeQ8bX3LwCV+F81YoTnTF
U4exDsIjeO51BUUWLfdBXYW5e5ssq4X4duLnLUNCZG5vodxSDEIFDVWZKdnxQcoyIvsN2D/sSrCq
FRIrZHLaIisOo+72Oc6wYGal09K01PZOU85uGEuSA4gaUpDWa5nx8KlwIA7tMRCs0aMI8N3GVXXa
L9ptB7anD3TjDotSykE0BL0lK4zar5pm0uUcYG31m+BUDOHK0BAE73Y8ePrYmInxq8tHfbR7m8r2
o4t22Mxf+aoSbD0SVRyJ/PkKG5rD96uRQXpg1ZrDHBXbQL5Tj0rS5iuAP/4SMuRE7xKU0PzX4Bud
nf0yPBurl3tjJ3tTYBr9rnxyRMOxt+xGe7JKopPhSXOFliZXV5kdFi6hccEdoKKmt6VJVO9l/Cvi
3tq+usRkewAWY0qHrJrZluVvS7j8MVSemFUZv+mEemZuCpe8wGnZlB20ZCXdx3V6ktLZwlzVKdzS
KndZ+wBDkCvDVfzTlgwOBS7PvipJ60aMDwfJmuHntECCmsUrzXbdsJqqbNgQ15SIZ02hDkgIDsSW
f7c/zAIsMNM/ofRvZdtYPn18cI6qC4+I5eCoSHQ5GosAauYQx6zr9swQXlLGZUGoU8jdcsF9y++d
JBl/X52sfBmC1my14+uKcOhzDtji1z7VKQ0/vTL/jiQtOCMpTeroG9xhRoLVxFXogRhicEXvitMY
kNGfuAMgDzQZhOclg2HKtZXFTw9wt/ozNG40jXvIBnEEu1KxrsrxMROshbh294y4G9Kezt3un55l
uAJf05q+eXDMZmr1whq6pRN48aaAvLsSfPjnadv9J8V4Jwj1pCG2lz9sMVFsHAJTk3NG7LktPL8v
f4kPN1cAHAHzTBj7q+MiO+z6H445CrrdlSC5/0i9RSILXdC3xZtowzrjteQnz8aDDiBfiN44VPe5
PhBH+fB2TgLs9U4+nsp7vvUKDxrQA7hnlG/WH+08j+Ae7rRVBwUITvUHrROkBGis5Hmiq48016qb
cbpWPuXJFKQrp1l1JxxDagtnt3QrzrZ/2GM7EhB9/C2a4ZeWn6IlfYPk/0RNdpN9jt/+VqkiXSpJ
tm7ZTvz9oGYDMmGFm4tIdTiPu6Ic+cVP0r0q5IbWy6Glha4EmExhGFYU2bHKcK3/ULQV/SZnqYcK
e8pLJnrfu19gvWfBWUQdm32kuOyMdMbh/zH0c83vAINbGtT3pSxAjmC20735w9zfDKPibo45eNsA
aqI3Zkdi++IcpmbJKDIdxIOHCnRICuaiT3yhbCZJtx4wp4wy1/FVRMgYpZ//6AcwPQ7rJZib/yBa
6zpDXTI24f3HZ/ZskC2oRtWHWWfP9hbjBbsO57GkNgvyxjsj5a4jtUZiltHMmfYYtnc+uHZTV8oi
E0qDQRf0nVLptcM74xakUpA25D/oa8r6ryEDAei8E7YigdUb8pTx0phbWHh6LE3EXyNOEdt8g06I
siIcgHyQunq7WmaLaA0CzGLx6bb3cHEexgHqw+lSP/6bq1fmK/MDAYSu5saTbAY8KmrGfCSFD1F8
QKzrsAQK+ppYuwVooKbzXlKMNAtW+4Gd2j4HxcsV7Tu5ET3+AtFHZv2jehR0MGi1ACzZbj7DEpM5
5owWhkIiYeVPCsmU0/URU7+zERq7hpds0HzmKsD9dweajX3aMv9JrpCDkm+EZBiiTEOJQQtWVbAc
i7TWDU48V+k9IbHDnG/nlrgCBhIAbGEnNLb2CDIR/yN9iAR2qpkglWo7d3DVyJ0ECa3WrClPOEfh
ut+gYv1iI5mHcmznWXEsDP5fIicqOvpLCkY4+44LnsLPYQTJ7rls4Wuc8xgJLP1VGxPKAO+O13wz
GBYn8fNYzMxJnM2pUKP+Xwtxx2aYerqa+ogtdOemiCLNpwqW6eeV1oIgVe8aucjaTy/+3ItRyblc
BI2SXD6MlqpidAIuiGR5MyM03xfy94beha97caoqtALwz1S31GTh9Kb0ByUghg0OiRdcQWmkP+c3
Ufv2U+Wp4/dDs7fRtjCT+gqI/NA4Y8qc433OSG1Ufa6ABgW4f3OG0SlCMFfT6ebV7rr43qptrbAz
9w7pcXfUF1tlOHk4Da3LT+n7cQlHXqbEV+tJSPjjEOpvKwBaATM8UHI9f/Ecy90tih8xt6d5F8rL
FQ9GBrvNIENn8X2OMjkqqN4L/+34/pzISEq8adas65LjiE/R78V9CHh7h/rTS+/krS78w9gsLNZf
5onk647mi3MCdc4I3K1lj12JGMp3fpmF/pRMKqlLKKFrmz99Oh7iumqjLavXczmh64DRurrvZ+YP
4C+i+pZUWhNpapiPh7t0DMJXlNcyQ7INxSlUD8W8svLhosz2Jj9hasSrANrXGuX25tfO6vIfjzBO
DNV/sje4TQ9jEcLLIPyuD1WqV0Z7F9MOvXN64Q5/ipgNNbjQgOEDw8ITWx5fU+xKbBDOaLotGLsP
fq8ncCE5iX59hUOm4Hzt5DrPIquTXttXsDMT3gdtEwmKtZcYAmrCUYO5sDwgmxmbpslhuMQzHP5m
vWBFbx8k3eaD0mh+TPBZd0bIopUIGALLyWac93kuDNhJNCqpkwqLoqwftLL7AaDNUvLxajJar/sS
Ymb0jai22WwUTrpH+SyC8DRIjsRXlM/zcEkDdhiE4SxdA9XiZQQJjsrrz1JydCFX9XqAbMRfvlyR
qjH5mj67pLt2d5sZ7gzb6nXV5U6IjDLTS2JdK7g0ThALeSiuMMeUmJDTR0DyUSJxwhMEZ5VazvcW
G+l2nAa5VlzpCwux9FU139gRlAE7cTJ6pxa4UqU/AemdY++XdTYbjMFURoy1SRQz4PU2OAng5Soj
mp/AIWBMJD0t0/RJXHkh9s8vuFMAiCWJMFwTuB0PSB0TIMfWq2I5N36ayzCUBFy0zgrdaZKEozB/
m3NI6WgVzfxj/E+2zvG7jvxX72UYz53ky6SkBZceUFKPx9slDw9aua3INxLdeguY412Ng0OHTCD7
afmlhXl/D7PeqECw68EazzEoHMVOcZJ42+ZAVzJVQ5eMcB0UDmgD6Npy8HKrvo3ElOXt/anQEysF
5RMMQ05Ps0LbG9ALKLbbLF5+FtLtEN23mtjaIL+6poWnJHKRPC5nBy68myJUfpNHwHmadTbMcbXq
VsWo7dc2eEzJLPFo17DKAi4fHdjIaUQuu7aG+UjrrGJYtlSXYfVxeAlZ/HaJzeGMM///vHB0LWIS
locK+rkVCuI5Yw/y9TmvvPGZUvYwpvgQMjpTE1/A/yahHO44YVFZ/F7atvYBNBsf9GI7nP5hTFTp
ENK/svRV1yeBEgBxNB0QFn45OfZ125ubLyY0tu55e30s2Ec9uzy/PLsDFJRq7MLeFMhiBHPYkadl
BBk/xOwcMG89xUgts+aUboF0kiy0JZP9UEf5Mu16JcbAT/lxyXeM/KWqaRIjMfbdGBkWwB2TH9AL
6Nu/f9SHygXYqQmqRXz/iYk99Y986BTlKeb2XjqPJYmLawwUXha9EaiRyJa5nGymawLDcvSEmePN
JQLTRnYvupg2SIKquTdGU6b2c09UNBSFSCdKxpWeniRnEOd0PJDMZL+xLixMlHNJUW70owN75HLv
ORT8qF7Oe28DhwL6SJI3DD+HkXQk7oxkb3sss7BrNj4h5g0pYeXz85PEt+XqBhTdPkfi3cqRrdNz
EkbaPDzlV+GzzalxkFnWoJAi7VUGS5VXHyowG+uqBtZgosWIaBJzhVlm7buIqKYXBUb2FmZ9Qf+R
sEM102h1P07MWQUBh0FAREvCbqRlkWVSewAXXL/yf02P4wLtvVaS/ZxZzaUO6ZAdwHvRZnaa3OPo
eZHtm2TMpOuH4OlN4M1ZiChr1i4g/jy97rvhjrDawnVCSTSE1dnrH5rmz2Jc70MMihQr3F0bxJa5
4m+ig2OC5dGzxI5iyVb2VdZ1iwts6RdvTu8IcotY0+TlFdaTefcuRXPRRkbf42twvCGlQ+DyciA8
jUEXyx3kyMZMuzKT3eyKWQyV4xEqOlTAoEXEFKM0U7I8rwZVkObFJHol5yESmEdemWRbup8nKvM8
+O40pAl49JVUzo/tWfZt3qYnzCuJK/x8GDbYA7oZctBFHGYRVMWOwi+4/Lok1AqpsSUgjmlabec/
R7Oh05nnJ+Tf3KtE2yZV7iAmudA2h7kb2C+8m9f160QM7nnMkkg26zdMUbj0EhR/FBMEEvYwW12/
vO87dMDdA+4nSsvUcwoik/yVJPSncqacsQfhz+RpwFWfaHk0EDg0z/FvFncKqr83zTMuLslO7CaC
0Sh0I3TxQrz63Qm0d8IuxvL9XXT9YpRfzg0zFnvSC7LcrfnKezHNhiWbcwo0OHhGfckPaucR1XDx
dU2JD1pkcRK4lcGAKUkSaxaYlZhVXNkqO14Rf3y7MIVrjpHxNpD1JYmo5KKiwToscwVMTrPcNByB
4pFuATFas3OZJxYAj4pr2ajlxCavyZQl6czt9kNsOriTdE72iL104R/NyBJu6vWZiqumeRR2w7Cj
UmCdurnmEkGhH59hWJLiUoqX5hiL0QjaSrIbB9AG+KhDP0K9tHNtIQdB3wVbSGO01TliPCS6UZEJ
bITCsMyMiRwxGFi49TD0NXRLsOMR6kDsCvdL9eaU4N72KFQw6rUcLNXg1hIqHNTXXWgTZfKYQJCX
lTFKLku6VyurYnTz0TT+Bzb6ymRVXNHgy6GaVrbSm2Uof+Z++trvRSYXl4KpktSVRiaTS/M+6REW
qAGBdl9GKgWxdtJu46Q0SVpQJqtGmZ3YrJg1/WRe1NX7JKgk9hvCUNLz9I64KMARVzvoJu+QGDGq
/x6vMDWUMPDiSb8z5kKv//OOLASPh20hHoUpUQE8Jt8DTB7Z6kDVadKuo2tsjtHzO9Mu9DzoxlSk
lgxn1SJRGX0KnlEYW3P+GsdxyzSUwZ9sKdo8awBjPRzRyCe5ukBsNq15ijJaTxrADwmLgqZcXf95
mxzcX6sMuy9mc9gN4uGx+WhApZ4EWsaPxG3RrfgWa/+tKKj4H8HRPsaaUKySgOZQVlnoe1TaSSWn
HgmafZ6i196chUzsHtpde+U/iHjwITvvQE5IC+S0gArmnQOP2tQfpU1mWzYm+WCrwAWYp9o4yR01
9S8h8m6kxL5CMggs4kXFikRhvvQpaDIhHa5L5UunhrsKGR/GZG8aZsQoScqZjdd/Mr0FlsHFkSvk
rBo0jOl+QE7UudfqheZQyznSIXEwyFW6sCcAlA0wWB2Upxmaa/dq4ARPBW6t74VVHAyh45D2JvL1
t94hIKEdcuxQRJeB693gEfT90zXvk0BV5a0wI2umxo4uMuSzcUod0GhPRE0CvP1vg33avaI0VcQY
EomPpNLuku2R2DaFQ3ePMRM2E/3TWjmh/buQt+OAIJmxpqQRVnABHFk3hDFGbrgL+VpoUakGnTKq
WjIcV2SlPjsxs9mYHedo7suBLWK48ZILD/xQjzgroV/JisU0a5dZHZzdvJYh4o+1+XMYEa/X8I2W
rf9dRusCx2zX/EV213PRFiRWwxPJSByyJ2u3pxxRnALxHgKQJH6LZX5Ch3BKfOOjgRhbzQqdgOri
/grHIGVopvvXwMHfqVtLwBaLBo0KUOf9fpvA9KIvfm/VKGNS2gXc8T8uDOMLqjvwwMFBKAeGeBcu
+HkzkfAIrdlNXoHnvqF6uoI9bNRHC3NZth5Nla+na7qUV7UP3h4TbSWGHXoY4vgwlnuJ0/KZogRE
hVv1VCDWW6makzjx/HJO5U1ohTuJ3eY20LrEMBY8Q4ogeLAiKGqTQa1EK2H6LkJK1AoPB1Rqa/5q
gI7hMkteaaA5rS9qhe+45TkQ2hbrPhbGbPj0a82P0J2vKNkoSR55PSAhMmSA4MTla409No0YzdGo
3OTH+6+jIIIjRaYZZoIGq9LR9VM6GxL80E3Puer3SEmb6XZ9swYIFZOaj3GEs5IqLqDq5nqTMGzc
FkNLDhFOP10bBPejYGw3EWbQJ7BE2o6/yc32wZfI8sgafIYgCNXwX4bbcbYWL1VcxTd39N6CccY3
2CXWf4KKLl7dhgtaU/tNpwLGgCbWIkKcoEmq5MNfRPaoufA8Xa8PyxGWbuOqUlsV3S37knzWk97t
u6pffJXnu63fGhoK5izFtylNkCkL4GziFuYHUNJKJeyOTB2XR1imQ8VSXMx7xbGX/o8Tca/5uPaQ
kONYjb33FX33HyiDS7F6De6PZlUpckw251W4RmfNckVl72fUm6D7gWvl599StrnsYVkwGgDYfkcb
B/ybc6EdGmbvjOSZXPkyV1JTDRTS4MwuKtjX3W94+CzHmG1dZ+Cs3PfNNGOt0qXCfj0lo5DicR2i
dFlE3bjqdq9TMxJT1FdBR/63AqNzHaHb8iefZ9XHnoF+Eic5f15BIa8Tv7d3O3Y9PKLhMELVpHdZ
hCmk6lRPghPqup5YpPT3yS9JzYonU7ihr9l5jqB5P74xtKhpgS3/c4byDUlgtX9N7yt4iq046fzg
Kd3/70zt5o1e6Jt2YGClIh7qv85Om8A6qK7lwBm2ynWXLu1iUIt/+svilusjzxnFqsvM4+mNCGNb
2o0T6UpkGf3QIO0d8EMzA0T0mFIKchIQwZbUcMzn15iTZqtIcTxVxw4Ucg5dyKdc8BDm/q8ehxAA
g85bPUE6Tf5XrS9CsAt4e/Y7mTEA6ROO0w5Cw1VkjSTlgrJPtDDsCG5Z2Du2KAYhnTDLYI1O/+22
7xOaKiLK458rhu61znleEmumzIkv1PnxfzHAZEmVDMkUTtYKDie3Ef4ygK/yCzeXJUoFwFvKjst3
n6gq/pJhe9MrzoZxCjlSaSeTo6nTKCCdCNoJrOdVw6DqCzUCMc6KUnHa3dBqT93PnTGO0thcxHDv
leWP/qFA/9o29FfiyLOrqPM18ObLrg2xJphibv39xuVtW13ZND9FrueW2Uu6aYVIeHK6odjQwxw9
2+Esr4pVN52uecZHKQga6QkO2MKFGdSvfa8uHAyCIa2NvCM1vDJ8rYVLXS4XvfhVML+/f/mVLlx4
PBDAOUL2v0xW9EDoJBhrIhAyo+lmgOQ9kYPSV+ypzOuuY/FOYo3xclA0gv3xFpoj0uISJbqJbBT+
K9qxhSIWbqyUbBf2ue6HoUNTmu/aW4kVbC9nvSaAbTLG/XsBWHSUVgVS21Pf5X7cIFtDcFORPsti
4+b9NYOusmMTenY2Mo9FBPRq8WcVueCSoC3FHUKEhDYGi4B4bNOdrrvpkhuPHLhc0uDaYxzW/oM+
mwFoLEt4wPupvOFzYEFon4cIz0YlAVNvTNTFG36JmIpaMyiez65Cm+VSr8tMSW5CcHs5Ckz6da7y
dDWEKXtd77AfgxJHSVhdZEpf8XfQ3oU21m5A/eQ/J3lFTGzhVDIMvAt0dr/gN6jLk6URYaKazBrS
F/vMFtuVVYCOVyU27RfyQ4kWKAig3A6h9tTpne4Q/ErgruCvcaEtQEvT8ANbZXy5CfFCLrzJAB3M
egE0MmLe/YLzKUpjOVSRIgue2csb/u2hRtSkgnFhDpq0HyXONVja8sNlrp7U2fJ13gWFRrMuHZKY
T9mxTD3N/MPcexi17g4fpKKVSAzcJo8RvUxnzNgM7tsFXq5cehOPAY+to7KRubiGxjqCnCHKwrVI
l84ecze+jsfMjtnnXDPvO6tXRorzOHsqEVgJOQfwV8ert6twCvvib9qcCDBy9ySwPeoXeLmYDRtC
kyCkCfxjmp6RYLuxvSez69gshjmAMCdtkvVfuWsrcNhRJs4Q68LpuBaeeXBQubkyWRaLqMIOCjjs
PHggaIuI+vRcDwELaerKdOoqOjFdmF6vDzlYIyTY68kjt/MLktGl1AxYOb2zcoC8MyMbqcLp/plJ
S//CbrhNQvA0ItA4Vy/W5l9H4we5xmNwKHQlLc32iL2bePVCmxNuR/nPv/QppQt+3nR3njyivha2
LysWFIoa96RLAoAWTnHJGJBR3XRZmWXm8jUof0iVWhKkEaiP3bdXYNieZNmQF3aHVp+Y2ZXZfW6I
oNCnlnFB0gE4zae30lXljp3FbayCCEN9C/b4/Ii5jPoJEmgr+shHoTAANLde4gZoh0XuofL9Ru3l
jKNHqV0YR58skZCnHqXd28T7mi6NdplnWjxUDzVHkP/jsaaydf/AJiBvyjv9VboFqy1PW80Fuucg
uOczDABbg9qQFqCx7WP3DYFpcPySN+gWQM2NnedrhzSBXbHkJkqHwpu53K47TAxnvRb5Mjcbr0mw
Lm3P7ZR4t+sF0r5WT56kiGbEs4se4WB7lOACcvFETrqv++O2BnWMBFJ59MfziRkBlHRCdtiR4c9/
JFmny5oQ+N/C1UgCisDQlrMKWNsRvnwB+jE5KiNF9MAeN/45nLnSiWhRZaezIVHHl1AQuldf8Kno
chCidAxX4UiqMC0njB4h2VhSBK9DsWV/vyJeQ0fOC7BZDHJWoyquVjdiTuUbk2AJv91KC2Slcume
22UkTqOqSL432DLrF/WCWf9v9ML2Qnf4F+u6PnNJkXqN5IdnAumJlZx7C9vgcNJ9LfQ2yxVHO+nd
K3UWes34cNvPgtv3/hhWr78U+QMtteKHppGg9JkYKd9Zg8xZRb5UULju2u+6CjQIpCA6zCvHUR+G
iquTDx/NjwleIk7JDR3NYCl7cB85bF+BgztmJh+LBQjZ9Zsa4XEtUeYcAHq7V1m1be7msvjASW7W
ysqaEbBidTgPKyV4txB7MpJ038EeGFSOMYuslp1KOq3OmHewY5T4HOFxImSQ8xTDpBb+Vct+HCpb
xjIElS3hgh1Fdu+fvZbplXxZ9x570QBYBPt1F8qGDwsE1W/Z7VLPTqUSDAJ0AXo6M7/Gb2u4XutJ
bI48/BIqlgFkWXx2RNHJp8YYQfPU2FC7G5lm8IimOzCguIDdznhNzt6yEunqO3UBDaL8Gdo7qU8B
1f//ybr4NcQ1F2jZlh2cIiB+wlVZzi0+yMl4Hi4+pAK5tpJNfk0/iQphtdhAkGqfgRE7FRy3332y
/Qv1S47s3fUOdPrX/GHgJJYEHQq+EZhZ2hyx8bLeJoEqrwuJm2E6tCywg6BFRo8E3Empp3fOfdrQ
PXT487ba78MhWEsUOp2R4RjAfc6hZY0JpSvb0D4upCqB+aqtQl+riMDrlPyEIs5JnuYXzvLIH9C4
9hqCmoc01lfDRdTrFsInOB0+BLO8K2vqk1z+gRq+/2RjIuNBHwAdCodFLVeR7Pc3IC6bGHJvPfgu
0w6Jy9DPBDxj0slOrpA/UVtWZb7t167x3pBhZ4z+yV3neFH/+wXC0RtCkoKMitCWhoN/eCkcyuHA
fr0UKnASHSCeBW+sFl8vt062aHO2xwDOT/S+b+x0SM6NmBvy0uX11XxRrPgKvN21YILWMRafFiGD
XsgpKLEh0yPaShc56dEHljOkYkMMsu6vqTw6ekssG73YQXnNwS+MWfdQknDxVTPTK4QKHrLA5vSl
8CLoefol4/3qzhn/ALco3/J2VKmesWnkHHUxlYUOEHAXszGJLhPl6kqsxcTv9Cq5DXIAx55VTICK
ajoCHyoAatJ4aP0gK31rPOHHoyLUJydcIQd0yZJDP/1va4ritRyu099DD9rCTNxQL+uM2gW8EfpP
t6PNO0DR5/nZRSeb56yhva4J2igahpxUpPwFXVe12V6P7/4t6da9sHoYa5JsM/SvmizQp9wvNqhE
PCNhL1QFbCmsYZlLTthTfHqDwPp5OtpCEWX4EqACvXxyohdkIPoYuyXnWaP0KlY+wuxsiaYNUcdi
qepinzDNJf7l+zVXDsaUw+qUFcdy0ZkMo+XyLUU7nzRbGs8QHWkKO8VC+pdJ/YwS+aupmFfQBIpX
x8ifOXVh+x9R3Jf7upXGE2qRjYg2og4aak3RD96HYyrRka6XkEs174kX9rJUqg5b67vTlIsL97lf
qBHl1yZDRbmG56fHKKmauxzUYnP3m3z1wD2lKNIB4apEXzXvjTSjI2yHYh7IUtSTK3V7tL581ioD
VUqISNsBqlhZnEJfsHmG0fONmp+ZTv4ugtYgHLYXzuT5PpXUo29WvITr2aMyv5bbwIBmZr0oS6cq
xN1zf+ouVwT/GP62KzARjFPilToe39xqPDGqZpLY6pkPXV456qJE5Ldy3UDfuwJAsIfAoFOasamg
xY42vF/W1H0+atiEJ2RVVciZ2qsKODsNlLT3BBPtkhIOdjoWxGFmBVbSVS61WMgaw6yTlCyPEXFC
59cSRcLqwKsbl1zNjiKSQf8v8rP+kGpjsmJg8vVBFnU2bJiRPXSoKEHPdOzJesFaLdqMCqibBZJR
2LXrM/mGLm6I3pOY69P/n/9JL83/6lNDpQG2svnUySY1UGt2HnMjWIvWHmX24/5kRwlwa/Fxjxow
iJwe91GuRtKskV4+ndMS/fU/qgd/xnvSWUpLEsX/+KiuO01TlaqLQiYJJ2SJAwKfvZWefWJ2JJjO
4mXcCSs2NzPeUcKkerQtNt5/sQvt15NmjskNcpXVnUcTYU7HUl6B0OdImHuyJPE2bsypQY7n/UsZ
AmlCHOTQZcQqjH/T0QwUe1ZI2F4pTKsFCZxusvGSCx/ZDOWUENCY9g0ReSrvvGTsX6nRwYL2TevP
c5Q2wlbgQrQLEa94ZYke0Vp1+EaVxn2QtWWKcBwI893UYSqRDuHnis+rCgSIIEgB2KdQq46KsDIt
ZpbF1IRw7mOh/eAI2TDXVq4Tag/51+L8pww2eHmgAOYYv13ehKiuOqh4M2RmEWb+nz6kW+CUZ5r+
bgUk+nc9prVvn6R4CFGm7iJIhBU3iw+u6u00JPoenIpoa8rH8kVrX0+zRPzyt5JkRsQCINoOI8PI
Kn3vI+QVRhyYMl6wDN6Iex8EHwb5jquXstIyiO7UKlUTkaCQDcX9aPmjtYBlsRwigsQcbySoH6I7
n1rgyAYKPnP6W3a0Q8DtNZkEOtoovA7JvvpI7ABp3vqCnZdIciwc1AQIPG+NFbliJUMIwxzRt7zW
/F96vTQfmLuO132vGLaumN61A7l6QkA+Hq/iFHXQOwjWqomcSSGjVwGVfsp9GKuFO3QIe+ub0XuV
tKWzKnNXKohvOhJQ6fYb6X/KPWwAKglDL5n6l7eI98CptaQmmoRz45XgVPUlK6IJpXC65u1Qvobk
2U9fVVuSpQPd0bHIV4E07eRltVBO/1FpxEcM/Us0ah79D/Okpg1ntj/aDXklYPWgP0TjnEo+rtio
xtPYBsP2mvcUGLCZMgpMfiOKcXKmuAn80UyhTK6akx0t2H1sfMOsmp0fiBEsAi56pWPlJy9+iKkz
Vq1+qtq12I063Uo+t56RZYfCzzXemCiaLJJ8k35eAanzbwcHCMD1UtkyM0dBv2rL8a50kaqgt8o1
3K539ZmOSrAMmdD6Get7BRUxF0QK+S/P92Mahn8cnq03PqkRYOn24bLSHlgQewhGqpt447BsXV6k
ifCpZwXzv+1JLzpSfwKYXgQigqF/RoNetcsMgZoBICSs0BphjI/2sY3Rt0qjGDhbhufftgqm9qaZ
hCHULyIqo+0SMq0zsJMEtgYfd3E+RPTe6znruWaAek5UUBPsJLo9OmhYIyop6omtnx9LB2H/ac4Z
U/6uvQJBAV4GNXva5gkIOle05Dt3mH7GeLkQRYRvNcYu+UViJQ0TdBVrKVOujgpYi4UsIfBo0A46
oZyvEtuvZZWBLrEIz/Qpu3hudbvYuHM3+TD4+OcIRmdcXO0ioLGWQG7VRsFHBSjQAucD1KGfL3CN
fUVDOf0LJxX1OKOzw2XGLDrw3o7D9JtcHu8MUc5dTTg4E5jeyif5JsCUwgoH7D14+9JJyIfPwKlh
6zFuLEPPKXdPuIsQuACkmlfGnInIrHYgCJUiM/hMvKyUGmqz/J9yKnEjdTFHtf8xLsxlycA0AUVl
DEY2XSPvtwQN5X29u0QcyhjC2iwUtqgR04Iy9MmeR3s5urQuaGcmo0ksfn8kc53cxlWBj13AlU5H
fJlouns+tEErJT+6wa950HasQw7ivcKv3hzhnjFuEr+/uMOjUmbcZ9/V/IE1RLpBkoweQ15Wd5gt
jAomYTnr1pHPgELB6TnW9F8X4k2byfQAPKkmdgBgWt2+tkfXa8J9Ph3X3QD5vkRNhamskH3BoyCM
S/Ic5MQcILg8KLkIhumEA0/hDGzAUTkkSg9HLDeFh5+6KoIq1CHitJ3GU2b2MK+CQa7n971ec/8j
z6EOQmrTmgsHYnuhP6mhhzvuBhQt6qIQe1gUrh9ZZg+pOZaS+pzLLkOjv1gSkGlHQWpHkLs7f1A8
uBC2NS2X8BRPk1FmdxdA9aTxyZnF/PLl+blmIEcovTC4ZT1M00ca1gtTHbllmBggYFBxmOzIS3aD
Bfhk3NHB4WDotMXxxUZyAsHoCmpKZohEQNkIhChMWlvlt7dbH8neUeQWWtOFj01RS0IW4JrNsApX
nmqC4HAe048qPTmqgNbjE3qZag8ArBtfrFOUAY75/ve4WRKKcISUEL4yLgTgVbIcJYDWbkZ8NR9f
eO5+xbga5K3K0ZfXFAtMstv10q9Zzi+jG4AaGR0pcRStLglpzNlUOgadHPDtlym461j59m1dYgSQ
fXwn8JxZ9F/X61WSoIyhMpPc31vi1wetkwwUA4IrlzN445qS3OMLSNGu1G2LENKEFNG1/stH1sQn
yWqSwInpOqx9qHhP+oYbuF3ELgYqNC/LBxMoGOjtMwDtjFfXVbJPLdyPVA4LvrNKEQqKd3HKe4s6
pbI/aaWLVp+i1Fuhb2vjqTGksjlZJzOHFVrr7jr0UHdOhUKRLPZBEtpMW6bY7t4qJmmXvSTL8alP
EONN4yeDzhSpg8+xYC92PMQjEISBUmIhs9fAxnVL2ZrnagT1UPwq81kD7rNX00u8M/HRLKGwZtTI
KEJ4i+bLCuD6rz9Zkly/Admu/aF2g1GhELnH8+ljIf93CC2G9TxCKQ9htbKG+E2jh8TLeE6pmBQv
3waobjdgP6/LxdgLUaDI2fKsRx5cbsJtBZelJuspDBXPPbe6f7VU42YJ2E31ZE0ryHSMqhFgpeT0
pG68f9EXIDh1oIjVDACYb324P9Aikq+aM8475yE9Bm39GWamQZrZCF3pYIpzKg2GDbDJLWulxc2m
JATtYZAGU/gfFCvYxq8N3nHJJwaELQ0bf6IWjHokH06jAOr9RLq53BvhBcHSQi6EMYQvZgZjz/aj
l0rGDrZETwP5Muv5Zx/sachasbUPNefnc1xAhYZmeDXMtXNdGdfIF4PK38ldd9XLiA69ynoRcxml
ZEaDoCjEcl1y8MkbCtAnGvihJ59GXCA+Gx1W14U7f09NFNWwyfEuxe/vVf9M1hgC75p07SRwPGqM
f8UnZw1l210DlqZD4yWjgw0t+6UCo8wimmMtDGTSp+xpYAZ1aDL6rSSFI/UmroU0afXwxbtuzWuZ
5irLw19wLU5zyRUkRO0ngzeQYKBhtAGDF1+Zm/78MeC59/gGJ/hsM1p3aEvtS38ryKUIdMK1yn0R
IZ2+7YX8hFDexK4FSFOEt8YlM6z3PBhdCNrotE8LUS36KkuHbm65BuEISNxKkrGK8Jpd87xLozxx
fK0CuphtJ9RaeOfHm8weT3JMapAW+UAK3HPgkvRKqlC/lClDGC9axX6OqHOjrswoWwfU93GB9KRK
9T+sKZtJydB2qfU/uvcJv2wV54RkfW6d1sjUULWEEzMUodxIQXzOD9/mEH+K9SXq8XrlOOIf7LqQ
zJi3cjNs3fdFoeJlRDkHRu5mslP1AVzBzYowiV2XIiDJIzB4S7OVGSiFxo2LeygTwHhBkA6V/8NV
adRYgPgGmqU9lAW4NwvxhL2eQuATxQvdtnopBwSADIm5wSa70QDSvFYtv2uRg0pJP7Tqk2ygDDBP
vzYFZkC0P/z2emwfhMnncn95w2JOH0gGUHjOtFGV4//hTAwHMKchVsXYO7AFejtWBh7KD17kq7kd
IYeWqW6Coso5/lr3LAM4sOC37z8yLeXOhFJEbFvVRM80EfokH4NwuH9KjXA3K7D919jjtNezA9+m
nYNwIqdPaYz6YckyU/wHZxKurEUPat2R/D22odb8vjZh7z7Y7KAIcNGZF0K07l1Xh3CRV7J143yf
rRSO+77KjKDRAoqYrKutjNIKqM2vNtGAmWkhfTRxSrsYVV5kMun0je56eIT/hqLrwoVn408IusyL
HIJOjMV8R9/AsSasoIUC/T2/LHf/rK6/UPzMu9kixCmwWhaJMlo2Ltqs7atBEJBNapzknIGUFzcN
CMImCQswRu37OfW5RcOiBsQxvjpZju1ZIsX1flJH8hVY/RaGnSRlMPNjieKM98pcFZkPGpMC2RBt
s1ieVDRoqaoENzy9cA6beqikGXRirbF2wedMuOvStDsA4FAXqWAmGdD4FZ2e97rtmJ0hoy3dI5xz
ldT9DIqMFDCLfbuGAyO9+ta/uUjaiX5kk17VKO4IovnlIN3s55y0BFmTsyvdh4uMHlEVxF29U9aJ
RH/gFgqUHkJ7SslXxZiuqt7K0KIFC64Xu3Xm8Jb2Fx0dB/S8rq7/ZJqKn861q0x0JOUKPTUHBHyu
/GLlZ6rAXMoGIXCr2g3LrCoBIuNW/f8TWc+GEeD28OqucY9DTANiFEckuB52rsqr8F9g8VtoQN5J
I5KiJ9TvRHrBv8I9LQCg71N+Clta5DsSK52k1/gbf6K+OzRiS8VNKQYscZCz3ga7cHCvaxgZs2Xp
r7t/2pJnIdC6ndM+vkuyTl80/hKYfiQ0ksvxmrTLifhTmx/q4RzzSPGGwFv9G3sQf53CjfDe51TM
6WeVFUUs33XSSXH+l7Jdp+z20TKeZB8AWFb+nOjXX/FcP1B+Y4Za2tGT1mSI+/svR9qjkcWl76vj
Dri4C0PIvmLNZUY4WL/cVm1pTG7CglQENRMKIiTM6W9bEmV1YVgXPlMyLxklMDpQCpVMy2hdd2D3
h6sraqWRGg9IbcPNkz7dVps5CvgnCp59k7Gn42llP0Hq9D1s/oJSIs+rAzQppZNg6tgSWM/rvHTC
CeuNoNMJw3K/A0kgF2Z8EdulZa7uDjjLpx0X7a1hOmFR4H2oV0Yb5XOfbxW0bf61ayek+GBsJ7Mv
edDb/lf1jWWE1VSi4DL4bciohBJvne7zRIyAZGqlsjrHX/URvYwdwPR0oi2STexzKKzorBKH+g4A
GCii+p7F20OBg2I7VEN3r7OP00dccZKIWJx3YPaGVyGbhIl93KFnBjl/Daqo6rJMHDs07YQrHb92
6us6PB6mii+2xjKF7UeyVMZHAXcnP3enlOqE9GLtT+waOgXvMlZF8ZyKDKjvJdubEY0gnYoWT82L
cZdB48gC1urEAjK50jq7AB0xKVAM7Keuy761DxXUEiOe5bhjk9zA9dlPvR0TlvmxaGLzmtGHXvUF
Ze7YaQ1tfaj5nVCigG6mI5oB3u8JPbsr6PVPVC6gL40sCNRkQqAirmgMw5s/SIxril7pJURcH9YT
7R2OvimgYxKotkV1quCOVIT/ikdnOiG7ViNGGKEEJi3C0ombgp0QkLAlyXgvKQ3jW8RyvmgRT/Lb
DBv73ISsiemPPU4UG6lASsjb8w1mQPRIDMc0UllYrxtcvaVqbkgaAhnSkgbogElyF00qTL1YdK/Z
ng0CDAoEvnxTkeeVxDXud1RyRZdof+cm/8fFuneWqe7BZAN4Je5rgAbyE2zM99QdNyEFt6DFs3hy
wXTKkgOpwKsBkiivKwzv/jTJ8doRTisKVcsHfZA0D94V9V9wUkWyYqJQorRO7a5rJztmrEgHu1zG
8xEEIEEAN8rju+VAbEitay3jxoOxTDFmfR3nCvAa8DHFyne8804C1CeiAyY7wk/NAUYW+eBvh+p2
H7YIzeFyNgJygB1i6IVq3q/8kHIofgaLz2LyatPd84urLj21z5r3/Si1uJ4MSGNNXj8br5TLEUPT
Wry650Kfux8J12IjbYaVUel2CY02WH8CREz3MSFZrd/x7KF5l+ivlWD8UZ6ZPY47/fgmXRE2HT4p
qGhwTtGV5DugQIIw/6t2fi8R9CaS5X155bmTel1UOPXqMAIx1Yq0s4LFpLfKVH/EF/th94SFe6mO
1G/t6HTcoR9B9owK+hyCBxOK6IFaSNqoq2a9/z32Do/kty8XqRsoOY/AbYNKb9q1S4H+2q7Eufda
fNcu8rmjOxC7u/oCuIdBecUk9I2lhHgwQPEm9r2YK8WyJZWskScmxDiNsQGnkab7YA4DRFMIQ5Lk
c0A/gQmtdI63TVz4x/ukSfgEQhRNINZMVaB208OtKAvtpojkLV3InAgSyOp/ifgUq/Gs3OgLPdUG
NH3OJ11nO0/BoinFqIy3tT9VmxINb2j9mk/TrwkztyjuIkZ8Kt31O+MtlI2DYTajjXzr6E6hiqs6
/YzmVZ+iQL8LqUoK/nmM+XxfvGG6wwIX/X1EOj7EBsf+kLiE0kP3KA5RMZ/BHFf7EjX6GC582sEy
MpsJ89nkH6J2zjDK+/XytpyUKblnGni5HuSHE9XIYKsbnX4PhGrHVW60CuTNqTAPyNXnwWMc4rKI
TLia2zPZx3gnV6TyhKNTZiO8pt/u1m06sgfQEaLiMUhQLSUuQFg/Hddt516eepVOqJdKSOZp5/tb
xF23NsGnWoZC9cS5VK/NKyefEB8tELTnSe8IgTGaXAaKZgqe/IXABl/ebBySKMNF7dq/CaHuZu5w
jKX2UTxeNakL+XRCj6wKGWWaybym1QtTLqMMMGQ8SUU4ruZ4MWnepU3PHGNG02ZMvD3jynIvUPqQ
xKxI6BsAbggD+WyBTu5y9v0SDFGN5ifF9vwtjlXQdSfdeU0mgHNDqN1oJaxp/86rCxYOcxIisRa6
xuH39ILbmaSvWnuzkhaFxc3ABqXJmXbloTst4a9heKWBB2muETbYFIrGFc1A21KmvA4enODYDnw+
LX4/ht6BS8j4hOCgV5Mf85yPYCnsxfo1uE0n14ojRcDGKDJyKi1AEJFJWJSoO6lACuQpFSqQgL6M
fgp40t0Sa4bKrVWSzIL7uG7GcgIAm0U7Ur/f2g/jYEPANJH64I42MxWQ2eMnyuRJVFG98viS4I/t
SSFtuPPDS/Z0pgLKIWlfqQCJEIO+63BhDVjO+ZLRi7GQnArzqfihKcD2ROZX/EFZrGa70uOVLz7w
z7PH6L1zX6KIwtoUeW2ViyGxjbpSpHURpZ/jslly5YT3hWHbXPmfTsGF4Ehkvoszr/lG5nD/i0gf
jsHc7fzaXFiGFj7O0QZNVo0Q/bkfV7p8G822qmP2BF4Ihx+fHMZdpurdnxLykndVVcDDnCaGfQdv
hkFu/+V51XkcWRsSMZbyPz8nhPIscY6wdoOuIYQ4qo4yXE7cpTv7pYSnhFZSM7b60HWY8Smq+mH/
yK3B7K9ZhAD5kV78iJA0XSL8HGgte+9d7gdTM7L0omz/1FAeGOxrI6j0SvtSZuq5ug0i/p+a20Mw
4U7u0q6l8ImxxFejwuQPEpUKaqkc0SVq7CNc3mHe92r375/158S/UOKEtNcYiqn4AoxZPjl1RoTA
RS9avdX2lcDNhVMM1LTXUKShYtXdAzygvHhAUJApa5g4zu0fBN1qIY1M4qngiPa+74Xs/mzrBg2f
PByXSZbdrMzrbiv46o02Nn7R+kAAmDh8lZCGic5G3aSPogtCHIMyccFhC1iOutS+JXRxRWXthISI
exelRYmsG0bU2e1S9/pgcZ78oE0G7SWzt0IvjCkuOhcD3gLbXb7CwnZlBZ1Hb0mMgbMdzJSgBLTu
HNdZ56Y8uRUu9REb67WCRJsyyVcGvQEfbFcWu37gFpm5oSDWEvLaW/cKNR/C63dew3ufdC/jIHus
WB5PylIIyGNRo3gLyOKG5hCySk/KyiwKdBEEEVC3GCFDsRHb/CQilVcT52bcdPY3SUzWTj7L2920
OWOImluvXDBtc1hY867RSJkDCz9lIYJHiXaimUBWu+owsIobzjQSZrX1nIEYFQHnUkD/YsRXPG85
rbsYaPiZeoSuEWdl1PkmAxoagIrKKIApGjtX0fxXJQSv98wNEeRgATMhT2QiVH0ZbvhU3A4kKH3m
k4DEExlEfKzmCFIKp5RWt48gtIxqr4zwGsO5euubKXmiZdKQcT/OwR6cILqv35L32XaqE2HwYuFk
lS8ll+HzJPYXD2YjPyRzu9Al4cdwig28nDAf3ztmaCzXivQl6Mn800/XEkuVOtcqHhNVZ86LQwdr
BZYgdi9d7lu1c4aPpF9MirN5mZuvmx5LZtkwecpeediThzV5DK/eA/Knx3r5wPp4pJKbDDGXwpc6
VG1rs5gJaHpWfjO+/1vP4DKxvYk5VkLlNuRLUhSSe+fOtw5rBOPVdC2N0vuZjzyMq8CZS83O65ty
6j247AU+S3ZBwMkohyh/BAyliWoWdK6uaSygGBv/9vMmvjsJ+F29REVr+cISmjzBQuMLk8iWyTOt
c20rGdMkEfg/awDcgMIdLUIqdbg46+H/g4Ka+RVweLXkW6yLvKRywKdC2C2Q7xAnVhtYNYZejDxY
glGAunjI2I21uMFzgKBqp8golOIqqQybAFsFtRJHYjqn8TrXg29kB41QdD7FEEI04vMgfIAH9/nP
kEwNjPABiE3c7xzQwqUaO1sjMChs5oxC7KJmzsV2/X4FQyDhZQZqpx9+B1CuI/8YS+FOCY+3GedN
bMg4YB0xsnDTp5Gg0hbjH70eswU1YNTuk5CREKAJYvYTGnDPYLmYQpGt0bmOYudbdRb08UwFIm5C
vAOp0mR+2MtNFYPHO1hcKqOgFcJOa2HOsJuHVXwe01FFv0g3NiHqbW0zDCwUqWE2nfdfzyIAdW6h
/rUn6q5uvrCcXOBu1lfcWNUGn1ZmI6yBLoIXw92JkquP8i3at5Hcp6DdZV7djfy6T6zqgep6l53r
l37ggcWOcYj9VBfFmdd+S3UkyR8LFIu1erDFEn1MLmguizFbNrFW7cyvvpcrCKGVg46mSojfCZqY
T0S01msTWQ+ikNxl3EjFKMZPBJzXJfX2KeVEXg9Sy3ha983XtIqM8v6u4rNAQFAxl15l8seql0k/
e9gulLQrywORbhVHmH1wL1DTX3O+TC3kh3J80IsdKLFBRaxTBFfd2prtN3a3ezDOhHgXRRpkIHh7
wGocEJzOz4CzCzPVXLGhkqMDGvP2f4srnwxdzW6rFCAD0jyLO+KHl1W61c1d/01gTDLdnNj8/ZVu
/FnCoUPzs4FWSrc8M7wxC61p6taRTga7pxbq1C9jrxAC4NN60VwYLS+bfQRR+LQ3afJlGHeg97rX
Wowfb4tk7jK7+BFRRkqUMc4ZZ8fB5D4V0wWE8ayFWnN43+yQHWGY5YyHgA42CUGStmDIDsiUrQ+C
GUlUzOAaDI+dyPFJ/qG0XnJ5QnJ7g4mt/qPoYfeG6YWqyO7ttUuYRpijuz2Qeddzh0PtDHADv1Nh
z6VGb+ujoONs7iYKsZGkf1CagDedazVEvlfShw7huu00ZhSo5IHk1KcbvhJZgNFGggKKwyFvQOBp
XMisJOhKcaEaWXMcuRMk6b8pYk3VbRIJ6Losw363etXpdJa4ZfaHYtqH4E5KngJR2t8PPyWfnhUP
hlaqN72gc8rapVhAPllWYiUWGPk9W/1PYn92ijC9sgdzcJei0Zqy+ue1UPQ5pb2O/gvOQWow+D3W
vxF45UHMvfxBjxivnFmrKSllyuDteMTa+r7FvGW8bHOCpR9S99D6in5I/g5h+lx9ugNLHfJXEpKU
bxWf7yZzzTbd5Z3PxVyJN4qdg8x5vRlO1L4LE4v3oxBx89L6qliZracIHIyHXis1ppYCzKdycVtN
myfS70kKoRArDiQ3G9Ol927sfT0mdKK6wTYN10h/pMsoqob5Hsr8uo4x2LSx709OTQFchlYH5Fle
zKVdnVaikyM18CkOVBL1rFkegrzt1ODNlC5Zt3tD2S9+A3o0bkPkgM3w5sk05NCRZoDGmDR7MGLd
iX5s8gR6f476RCpdmt/9X7h2wSm1XEM6TAHQnL3TapLIE1kicDdMs9/k2TfgWX3wVzKN+YTvwLtY
4wc2H+jBxFLtuT2Zmjg5EXc7g3HwpmH8meV9hJHXGyxm/mRtbWW7rqUtPtd/YF4gR0I1Ns9XfAtk
TidRIf4E2/FS6aUXkQEl5kMZO9K7SNJ66E9AmXMemTzdudB7O3sxrL1eF5ftl1ZKRd/ZUF4v3OFG
LHSPOKTxIt1fxXYfJEAQ8g9QLM9+rVtzVWSBOJLxwmZ6bJ8XZM3LE2uID33tOP+Qxs3KkXSbpX9r
RXEr76f+V5Q+X5ifyoR+qC0LN52bg+sKTtMJl89m+23VenDASTVB/262HnjfyhTFhVob9hQwGTzT
/5ke8H9PyFkY9dSGadZIDePtF2e2GKS+rjuwl2xoDV7LXiJSzeTFTbZH3jLN0NWxhddzX5eTOItS
2DF/+00YoRiqmxwtsBMUDpzwWiBWcLUL1hmfS1kvJyePS/W5gV00YnxI3q7OOW3uWqzw5c32P+c6
vbumDyjzNDW/XT5odD8Mtopk9UB9ohLQUJAkyXqV0RHh8e08R+xdJbes/8GWl6TAHkIGeoKjZef5
3LCYjuGbWaSQH7DU8QVvMWAOvx+eca4neK0WELAsGYZruyxI3ZaeY8NN/lU2mTZJm38EmgVNxME9
l7CYv+8iDJWMmbvMGz/bYEH3ont7oHWdzYC2qEOoIF6XKr4HFhjlaYoVbLQlqGrDIK05pEwEcVW1
7KkS7zcagHF2TNj855noV6zyNAxZzk3GAllTRMB71uVxJfLTJEmm3tXjazKN2/godGpB/oOPtv1p
r+ETmiV88EhbPf+Wx8nalCLWyv1wHq4DxR9CLtj+3c1wVEe0rcwNs/PCyBdCyCDbjcFFpRTjhnEw
9Cd+LHj0Y3OPbn5nTjhmaVT3554Fclr3SSzrHfPHnqOFJFwfLeGCzwq7B2nPV3p8I0dLytvMFFKo
mfr9Ml052xzEVq1OozyHRGUlxxaYmkH/dXWyZn/hH5+6qPjBLHHAVQb2XJT5ybQu3ZM6GBvDl7Ej
6BkNNBl2O4JnwQTkDTrV4qfpK7324nDFVSJOccYjgJtupNoMyaE/6MroubkSRyj0mWLulF3WoQmW
ot5ASKEpGP46+QVd/uNGgnCuZ9KL9fV3jjZs7qnySvPFpPonzDKMaQHYjOZaBxWzDJ+sj+m5KK3z
jilunQtiGoPYxvZwFfeQa6rgn0mFa6OXX8wWDa5x359IwstYqNwKEGH0dA7zWUarTW22/jSoC03c
rrR64YkE0morBKY2i2trSGlbhPwvtaB/aFxnACTAESgp0uGXMMgJ5rqzQUwHbS3us6wymMgmU6dw
E16EQsvl6XE2CQwLvobgX950TrLhfcZSGyJEUA83SZwRbkmYMasAn/xBZWS2Rwi9tIcHGcgYfm3O
3OkmYohguepisp/rhjPxoCN5hyHLF97h87KBL/sUQ0b/bP1PunkvmUQKJ2m/NWF1Ti/xfYaRtMnk
lfwdNIJappOHP5ez6lnMEkaGCPf/27TjTuirFSLaa6lxpGSF5Ab6CWEAHj/BoSqvzfVxXhzIwB4W
tV2XyAlz8OGjKa6b+DionPeW17hXZMuhy52JDY8isBOHlaLw5qu8GRiGZVHdWjlK3td2IlcTBIAl
YlvL5LFe75hRZfxQAXYwKco85KHN0FxPsHhRxtlaAdUnNrE636UUDz3ltCtIm3XZ6BOUy/7f6bIu
WzJzPhcE2p2O2aW6DVX26gw0OqDEk/DQ3lXbCMQfRwgyaLCMdvUixmv1UtFxY+g+sqVBzNc+nBdc
n4e885p32d/EvQCKoMzGxqGTjLKJMcuebuHfDarQbZdGJIskgndVvvLQDXPLyxgVX2PSqia2qMVb
BNbb50txMvVaLgKS7u1LI1oyrOKIg0cEHFr3KbZWkzyIUSOdLIu9fWm3+QSwF0DBkOt4SDyxGFuz
qy3kRSNGQw8qHFP9VcVe40QGxalV78Q8/8ONd8DK4T3+buE03YeaBJ+P1M9XXnYN7buJkK/kzlap
HAUzPiZbLHhQXBZAER6sa+w9DTLWpz8WS6Cs0Sl5FiMbDuwHrSKQTE9wf7aQaIuGwMyd4FU+yRZ1
U9ph/HqpCH+ZNK+ex1s87I4tGivZEMT2q5BmybOCAkycDj3fhnC9I5p8zU5QZXAYrcl9WEK0O7av
+xmFn/OZhIlYeexmCTZ5VQJ5Bbz8sLCm8TPDEyrx5rYKK1ZB64j1zosJCzth0jH3TsS9PW6Nlvz/
9vtbxrJS8il4pqQFn7HH9Q92Wrs2OXHlI08MprP+6c6S92+FcV55sXzfljWVb0eQL0Q1Do59jtXR
7KXQ0omT+vScHi3ezUmY8WucYASU8LDgip0je3R6vw4p3adLVHgae4BVsMT/CJxoTTpS/ukPkkqN
nbi7W/fAVZFF7MV5Z0OLfLgTZeQ3zeXvxs4c+6xd5oLjlvnKOppAIslt8H/ao4+JqSUo1kJHm4UI
d88WOXvMSITqBHYYjIkSYRqHvH5hRXXyjrCL30EPxNdJK3HzyvBKJgasSYpN6mYFAr3UBThYQzd/
VZiurSg6LppZGfo4aUHl48cFqW+Zxc1sRAzJWawL/FUiN5Z84g+t9IHSMkO5rGgZ1K9lVSxIlAB4
C7m5d+WoE4FYcc2cMVqI1pKRYDlt0m2FAIXGIupGh8RHEoxNKPxrMp1CTdMWG8xiUf5TnlBTjtao
3qRrmm14REJvnEZTccYzb7KRKRw9j50BP8fSpw6429wdM8RJo8Q87PIyqGQYpNnEId/xfbwOuQ5E
huYnLlZjX6xLY8k3STgurswj8/9kRBNbu/WBChKzleKjkGGeQxJzfdmy0zM9pHQXC5azTfJfzVDp
oKlWezlnNuvUGYa4eL7lX+an+KOZxrxrp7gdf47LXl/fiAl9L3Gde5Z/SRXpOOB/84ubf83oLdUm
mXuI1RVEseT2RcdGE5FbhSXlTPOadC3uVLxITPjBXAmTOAmzDZyOXCOovZTTER2PMbS19ihEhOg2
9Tovez1Id0q2f/HutngDoxApOMOibuDCRp1bv0nRmN/rj00LCfLtQZYXPLnfc5Ib+pHzShbhtwYV
PrVbknIzn8pkqdAY07bmi7Wk6MAt0D7LvOWqfxOELNJvatBwnCIM7B5yN4UbwLfVtJDOX0yE17iK
s1mJWgbLmraS7UhgbXRz4azMihincWbxRoWDyuEiCIhfWUAQrezTygqhIurEaXdnjTlL7PBihLaA
0WNfvQcsUmcoHQHi/rZG1IrxAOLjlehFIjynfNYDjCWJZNf2hJnGkZab43PhE0PeGkeKa3law63g
mCr/0WykXriGa2QUNmQZPkZayGZ9W0ZCEy061Yqx9RdYiMRot6ZfcEBw2kVKwhYHHgH8XcYXgBX5
1bzPtLCr4tONV6FyIPXjyCHCLbAE4biezTbG8Bu3Pq27xOO1QWLtgU9ongp5csjxbLyNRrY7F6oM
3bAtoPOEw9QeqQXpdeEahC4FUe6yivx/SAqVe48O6xtj+eu2/CjIjG5pfKwQnrRYPgnhxSqymEOY
0SzbefLBkuS0edjbnZ+Ut7LCOrm95VM0zBmKw8F3wGxgXNAcuG0ND1G6wx9ZyuSgza8ebXk9cf+a
Lsbzizbp0wYark0N15xNRtN0PnUuiC3NP3MDCJNeOXEde6WA44pO00i+F9LMTexokJyQJQIdu1AU
7JLr86ddpyFAAR034iJwlFuLa5v/YjYWOXJmWfxZIfJmJajcs0jeMmafU0+OQ188Ve7eDmyJ3ITe
Yft50nslnVo6LLqsSbzGUwNeKgDHl7Mcap3vzJJHwZQuJ8qL0Q+yxVgbJHE7wTQwiELXVoAsFoNt
wuX6ANad4Wfwqmz4Eu0Az5dQFEt3dQv0Br1i1UcE/YBkLWcJIwKpI9nOnbGnGRYDLGvZ/K4RtDLo
mBnuFF7kA15uf34iOJ0xuY4B8f61irrU4o1IOF5rP/KjgenCgFqClKzlbrRU4D6bduCF8ykH+V0+
kyWXv1PdnF7VVCYPR/ND/9pf+tK/yGpvdIACEDU52CpDUlmNlCFSPeczrrZoWl21AidD7a2TMmUY
VnS5HkHemKLeqOwO8+pQp/JOuh+WReznZV8MlDHO37yK+/FnFEqTNizijOQh/9/a83cH24qBmbww
uH4EtB0HzcXaSx1pQjTztQekx7ej694VJMRmAb9/8ebhfkmbr/JpcWyT3E/rkjsslyvQWXpHUIes
VJBfXEjOTiHoBlUoXGHKZ3oaQEJaZIUcbMkxe/v7C847Z3Uv5wFgeNl/8iCQo1z7sMMU1StePxmy
h3qMGZV0i5Yq28Srl22uUfAR9v/gzyynsMpgq9bhPoQThTCyu0DVFWONTQac+pS6/oTibD4Mu6xa
aIOzyVj2ndeOdIwSF5l9VpqPzuyo+ksL0vOG2pGeut9wDb8cSqFr1rmh/2Od4Jf0M3kdooN6eW0q
NX2+YRnMQTsFbB8ejoJndmKD35jRa1I/PJTGsaUFN0QA5hDyMEAc+fETMkXg/CreC56EU8WLmSOd
OLcoY9ZANLmgTvsWuH5wl0m6uLs2ztlAZXrP1bL+necqqgGmonVfxbgdr+RvaJbZi3GYiyFM5NJ2
V2sDxU11NLy32kktlO4hrUqplUyjgL7UgQSfAqbb9JorM55AG30b1Mu4KU9vC0I99j3yYSfI7X7U
OIRlyHxFGmuYFLE9LOLaNbjjPV/v6Wx7AGDUaaq6tT4XWpPa6xETGW2TkXNEHyUTltajaXjjjlDp
RKMnILklzCYVkQzQh9r1iaiH6lmRFL4cLCvYgVp54hRUHwe6yUFImHfMksrDB5OuQvxyiMV3lIJp
hTgev8XQO1gABSdbGp9Wje4i3wUwSA2wS2DG+DbJuWNxEoJnF/FlRvQdlBpj5Y7/NTR3D601Hf5P
l6I0y4o7PFmNzXUcpwwf3qYcrpthAC2KDp63XwffRpovm7cBg/ggOSY3cpuOR2mFl3eGAaJAv6lr
AopGhWVZf8L1L8m248wQ6BCK0PgGZ98Lr3bbeBrk6W7SBIguV0Y9IvrwGuShWebtpUUxfkOpVG/w
PA1RZAuh5KD3T9OoBefTBjcr3jEeAUsoBWnlwIYjyMuBRSWDLaNm5UYlOfQAmckvuBHzg2vjvfBT
02/fxrH+AXvIGjwtriQUVJMOLhx6YG39up9NN2XV7UrQiX+spguxEDzAvojyJfe9nUfimliD4K7o
k3GbMHoAyX88V5zcUl6fLaP9X+qq+nfYpyzg5oWxhAwa7j2pDoPO1s7CVpzHOfAKVvFIg7Y4oaSf
+gOOlgUsMr+sJJBAZxr6imwwpKxNmqEo7Q9QLujdBj600B1pWVX6pkmUElblB75n4SBD6WmNTn3r
+0TZZUsRL69y3FdmlUKpUI2ycTYLpwZNYdagHuWMcA2n5OSoT5dwxWN2q0342aTeG2yVFm8/FUNr
q/kIFqPhrQocm3192SrkbvlkhNOp1z3oapCJBS6Zz9Z/EKosyitdy6qLgPUoaM6adJmt9BgdxHMv
xCzVzkdF+RKWHG6die19Jvkh7x4AuRmsv9bL6JoD0xtjOpPL1/R/QHvyDB2V0c1ebeFZ27zWv6eF
D38MuOiYYNIQssdKk8ZQNeP5l8ADkKqBmXo7c+IHlLLk6NCJCZ54w97y5i4iBKZ+RL6m4ci265ay
XAJGgDUDDbbvXt9q2OBZ5BY1Fof46TwoX5Al4RJ3YUAUHbSbsneuSlY9T4dksmbGAzfaly5AoCzq
x0eKc+MGakhsWzULWdNTToEllDzZzyrR5hBr9DWsu7H354O4Q7Ejq1jDq5GrBrfz5mqB9oD1BcsE
4zZwfVr7tF1I/PoYI+dIUAxAcpzPgqeBA2XF6Tm5YilgJsFbMSF/9SIzyqIw3PjBpfuKMqwrw7NW
5OMsEyKDBVwVYXjSk8CnvHC4PEVX06C33VLSOKCT8HajU7eyvaJHlgqT+per4nssMZYQL3fh+dCg
H3Q/m+6oR1dCxpe0TkIxI6SclBSzSHFcY7mgLJkbxTuONneIydsK2SBERaxHXJFn7Ymfh0k5WVWe
NopNjPF0SzqhdnCzDLd6+Ler04j4pgMCTsfHkSRkdQmtpU1+ilq2Im7r7aA0hFz8yOb77NYxLKCt
yVCk6gr5ci7XdywYJqAWO2E03FGXT8c3H4iSDPSI05DSGMz8zjtQFHraUy9POIVnvUQem5btaA/u
+Zo88LBA6KuInyaqcrcMnPUopJsHGPZkSVXG2+XKdX3kWgTF8E5Hf2QvD7whwjAjkJIMvG9EfUcK
3NcXTqTvctK2/cqCutkIJyiFkXIGYh/Sz0CO+LV27ETWWxP1kUAH8VUKVKvXoftD1DczcoFbZWaF
fQ27ucEXP90yTfxK1ur5KKkuSKyVC2J8NEWgniBsUHCCXNf5dpF+UAuHJN5hViZYx9SEBYVS1Y1G
b4/ywznp0FeLQGJthmHgCUkTfVChxpNKwLbS/hr+pvQTHJ2rVJIEU0Ku2yqljnUdlykg/cxvQmhO
YX6GGoMAogVzQ9Cy4lA1gnSn6d55aMLcqbrVjZUqhwN8wqD3xHJD5ccFNpSnuamkd4H+Pr2Tyxwp
KHKXNxRhYXpUxIEF0OgSbchZSDdpuJIvkv9e0UvjThZ7Ef8FmzmCegwmBHSn+d0F237f1JbzPZHt
yScFC61TyVIQpzvdW+dvcB+4gJwhcEvIYPcBIGIx0tDM83qn4lr71SUkmWfZzJmQm7gMiRB8ikKz
tDErmhqVqYB8FLw4oitak2NkCi1XjifIq5qGESCJKe+mSTUpFrdVVozgAaGW8VPQsHL/g3wv4z/2
YEXFaiHHEyVvZwxobOvM0u89uzqvLN9LOg/rRd6g2XOiyG7s9r3IvNwu40jS9M1eAblgnEqV3X9d
l/7fvOh6FuH0BKWUDzl80o2O8Dqu0Eevjkhh9ElVnLPtbtBfzBpzhfsF8LouKcJvRIq8Vz1bIyz/
+SZuhONbJ8+imtZcf7+MVH6I8iA4spZIwtAB2BBw4VjPxcwFOjk1iaEhYg4B1ZbPSen0rFbP2CF1
Bitkja2Xa6HwAjM2QZnI5uyEG1E+KuHiNIyyZqYWVyvp2B6R2aoRXxCIrApNEi7eTKPhGs8uUFn1
XVjOk70NBegCMp5AVZgp6DFmu09NUp9q0ex+KSY55s8uLTpW9FXaLPEaXOTtrMUUCaUFmgtXe0Ey
dADgmOT0p8S4pKlGY/3Es2zZ2eZdBSO7pYWwyg0P5CI+vX2mkzlAUgiyHTk47dHCagmpyYf+D85f
gVhxRtg/jaYq+Jbh2yMXZsRxX/vwFdm/AGoNeF3NYjz4dN4wyklGFntYgXGNkARSLelArrSgdqf6
8ctSKX+xxDyhUbM5Ct91RVWuVUxX5VXSydUXtyruxTpirr5DudGwVw6R5cEaUl3ys5bcZ5wj9a45
Qg8Hmh9HLzYh1+bFMBYZVkd6Gte108928pd2swhsYDJliuUel8N0z47ChP/2NkhzffZapepcPYOJ
k6ubJfSVp3BfNMosyfUlt0SUUzf/39DO1t1lA1Py6/oevU5lwf6KSfejaPcsq5JQ+Wqk4HSvk8W+
jtrWx4xWYS1aOPFoUYpl1s/K0GUHlxh+CTeerw3e0NnRuBOTLwznV6DIaIhdS18s7KbIlzz6wV7v
wTkAbUC0X4B3LEgNGmqIDFzfYitoRJhorHdGqaFTqOZL5e0XG0DChASQRimnCtd2sMmyOI3ZtR+T
CL+FlAkhUtlLCcjUARjDARXtL+mSwbZqUgEAeKdo5rvLM8SJbRfV6RyRdJ2sqiYBAjnrXk2q09rK
sUQV7oPuxtVVYgXQ+/VLHfh1Bh7l4rEjfqSKn4bBC75pgCkfPFKcmSsJjzEsGA7F+i9uG+rUkQA0
c05qs+Wmgo2WNehw2fiFpXMyzPs7g3CH+tTQFQMsLJhtjADsSi4w7S07pBMtdwppeeJWnanC47/t
eU/OJNt2J5ZEzGojR2zyGLGI6/+hfjcLQJ+XEZgCK6B2wAVe9U1uObeRb3513W+ovPVjFxUT4fHX
IVz5B7cO8FlV/jeN0efWehvWYbnUPjvFQViAWTmGOmBbjZU4C6Vnwaro3Ml/a6oQtnUqtAMDZ7g1
jN8KH1vYILk6xlaXc58mAUKD3UCi43qJF+gHfJVHY6jI0Ng3dvKtVkoYFucBxlcpe8WGV7FXfuZ6
yUG0D0i5QjmaFfS7RBTxGhhub8L0j1Mr3soNly2W41NhiM83tG+LVjZSr7MJicLImQQCvsS2xqfJ
XjIQTdmbn1vxe3TDn8sgFjPDOsTTAATbFTl3aNgGuvBT59XDnmOOc8AijCYDWHaubl8adP/rVZMv
T0tBBXTtuoyK1OUiB/B/y61XtU/c1K82m2OkJJTO3zXbMGXd2LH1bFuaLQp028HjhO+1UG6oWfEJ
9dMfTr9RL1XwbZLoPYOykAgbJL1yputVb2silkWkkGBuBwyDYxlWXNUL0IBaYke00IvgXlk0eqMM
P++0ytcOiPh2C5BP98KF2CWuUyo+dMwZIHxX/g1yHHrvFicR1YhGwWayhEkuxiHBet6o6N+bAjHf
cG7LwZF/uUe1f00vdkImqJqZdZUufqd3baJHvAOwB3obwBghiaWbUa0luwMjDWVeyhk8BITrqyBr
Iz5lIu4FzPPLlMwHyHwPLt/wn/09thbIvDv5y02DpZyCGmShQGGQbzD1atPST8lkTxvUaQEbCfzD
2dO9X0ZgYblWpJ9xruJ285iAzL0OyD7KjxSlnGJodb/4RzswsfKpRGOdVZ7/lPJ3ftsN0c/p8Qp7
sKUySoueEnX9MM1MtxOr2dLsUR+L4PEv1I+1eyatRJpfdh2Iwk1ZUdhvADSHl0XqZG4cl0hGNrbb
0P3BJ3af0EvzPHnQDXpiW1PoFH4es5yGDipIE7haD+vHx/GsTsSHzCjMweZ21Bau39EOajCHVAMI
qPEqUlTWcjFDYVeQfI2dB7UMLz21cl7MUhIp2sEZ0tAhkGCaD/1USbU4Z66vaPvwNHViJTuFKlsK
7+XT54jARvv0XVRWCl8tc8E8iSVnAXqG53Y13ZZ5dxnx67qQkY/joTE7ga89OPueuFH668CRbEKa
i6S9E/fMCyFeqjndGshGa082LMWOc9b/j4h8HfIT6hrEPKqoMFEL+Gg1x9Zb0ZpvWnFPfSoLzVtS
oBgL9O51LR8fqZl811kwxRq7IQEWzsfoCthYq96qH+4QNsPFKnMmXnPWomXEb6KnkO79fr97ws/q
mV3iaH63ewGPDtHYry6Dol8C3Wtb3IWeJU/HfPdOwBbEIcaV+6HdCDXJMWNx3VxX1jO14mA5Q2DM
mo5BOmqxEei7qZmRrRzN7ZgQFKvP/7rD84HpVUHeNgRdXn73AskaiufHArr/v/KCNufSxAppUWF0
t4tuBRLPA16pMy/I1F3oRYTdspbll/VMrAdg8ZxO1mW9m8+md5gayXt04OhuzKiXBm4mt8pIZXyL
IVvixt1KS1oBbn7i3PX0Sf3HtklPAjAmRTBt6NpG5wo0wIrUKbGbtrhWQ7ClIBOQIh61Ohqile52
LJ96cfXf8D2yT3lBKCxXG1tSLit2k6celfzPUReWu2vx4bT4uRxWdfaBKZr3DwF6TqNc2Oj1YlAd
UB1z4HOwawSShZdX5gPxFXc5E+eXSi7wKpf8ADHMxopUE/SYJ27UTUrkUcxjIYn8Dvj4CHl3JhEH
k3rCaSHa5FV/mfN78A4SrAuOGHlXTtDfJUQlI9Gh7jaSFYh21j5HBvShfMF4ozrkLzYidvql3XvH
w33HOcp/arlpCvFeY20hh9LXiLCuOO92yq/jHv0iaybEfZYVN/6XHoufCI0rB4rwC3OORBmZJD0y
TVp1/WO+TrMH5oU4umNmdFfeF54saWMbEBtHqZt8dMFehUme5qN4IbtUrHUWGgZmG5cm2eG5P8xa
cGBt0yfTVgIltNSEFUF+egA5LLiQ5p7WoOavM6bIrOYpREPyUC+AW4IgS0sIR8mjOKDEQ2CiY951
9OUACrkfPgng4hQeVIfrTf73kCfeIMnK+tLHoAUSx856aGJpEQGSFkCLmy2iJBef4wuw/kMVlU7C
3miv1CqMOji3QDQFxrQrIMG78K8jdW8h7V7FmNWCapKNl2cTyQMVHcciFlEVaxAbvyP9g421kst9
MxGca85GRZCZckHRd8kEeabr6bTZ7jOc31nBTJdGR9HuP8M+xWsiL8YcZp0aBs+FH5G0YfCeEu2K
+Hky2rGe3ucNSABivWOzjInNnfhnB6AF5EzPS78rY4IGOTuE+WjRLSbfIuH2OppQPygbXfifpk0t
I7jzs7k9uXy5ZLtOQqaer7BETM9ZmtfFw4Woma5bYSowQ3maMXcksvTt9uot0tdC1YTykKFAgExR
UZFslNohkWiVdLBH0P6kXyEM472QdomMQJjTOJ8X4aLWGtGhPEwnBku6MFaP/txw7keXK0ucf68T
iSHCDQX1ADwEzg1H9/wPamEscZTJc4gcL3G33z4khwwX9gSAPcRJTbhdVMVjXPHs/8lWDFV9wcDc
TbvukvvQ/ba6D/F3QVoxEH4q0N3DyW+0LLnYkOk8RIYLHV0IVPay9nv5RjavC1uArv+HUoWA4JXI
U13dkuzMCFO59BZJBmi0Ufp/fP0j1FyevGJ1YW8OCzd9Clu89Cx4Drw0TxKHI5gP4W/vJpb8Gyf3
gLL7xlE/lpjqvU+5ABkuhAimpnyRVIah4VEkNDSqV+0hmrlmgtT8RLsrNesLYPglUzqgd7utxVdJ
UoJ2bbUGthoQ/macz8T3yQUVMaBhV8HKC9GkNekLiEwJWrknLdnh4SjiaGHZr7LDjppuIIMdpU22
ZI6e/aZNu1Isz/XsjHdN1Q3GOvbpOfDQC8SAdnMxS3ZszhAXJWjV0w5D4VnNeymCfy1lKjGZA6Tn
y7GCAAWsgFmbF0E9ZktXxXm+T+wbQtafidgPBETcGaSWPnxHSxxmgvKcDDFQzarAMTy6GIaroB8A
hexXiE+Af5oTfB1fl6WJkQcBbfm3WRGgILzfrm2Q7e+PonzlgJCIUwwS++Mu22pDorGB5ELinnTM
7Xbqn403BQ7Dfv84XGVYyk+1hlTm0EX7nocU8EfxhE4ok4odBZKZo/J4LhGci29uNJ5w7m6VBlXe
48JgESgoDq6iDCiwzcHOib9Vf8OvioEmeOLEKMSmsWUCKr/SEtdGfZrCFlLUKbfc/fqzWGO+R1Le
FAXMlqLrS4KIZTjD97rgu+UIyFfCyB9A1RxrF/4aHbDoK7gTBqQ40ApJhHnvD5Caf/Sitvp1UYLf
/EM6R7KrO2HP1UtaT52yGS4KjEUrWfHK1eeNJiDQZI6cU2bS8CXDiqmGrOm6sUxSZmTx2tXYomlG
w5n0DpNtvk/YDghkHX64k8LwoSuhYS4TEq5pe7ruPb8Z2eeOQlPevadQOmisg8jDEdXQh7R94MUH
ks31prxFYoCfiYxlE6pADi3febRA6eS+cLbEPtI3zyWpgTan6YkggwlLsKZ3IA8ibi8GSZW9Kw3E
BF+6XImK2afTyYylx/iemw9beu5hU+TF6hiluGATz5QBhgoWG7DuSwRLcM93M8jrttosM5RDk2r7
b8WiBjHZMC+jQVLOmGfiFlJKQlNme4sT6G/YnYYPHP25e1qcwYv5KTTqxdptj5lcqMoi8wEUK/SO
/w5PcsSUloAQ3+ujxp8X0mGig6HUmjA7Uf8LrwHwo1IAOU0UHB6lTxsrh1yxqHcEmI2UVa8M5sGH
5MtaFrjwTPK9DSJ9y0o/NA8/s+2Rn0xp69aBI/hWQGzkVFIUuZIbB6+uibXcwrErW7+xoZWXVodf
B2XOWow6irc1N8Avj4OWHV529aeTLSP8d9Ji7sJ2wD2vN7ysb/X8AncB5ixA9p7fEKwceqHCgtb/
mRwkI1YNC7cs6JYY151R1KMYPXvk1ior9MzYvESXk2PTWdbmbyE7SNYPU6cELYPRNS1lYNwrCEa+
0JtatFZNHdwHtBnEAeoloISbYVOCjKH5HaaEEamdjHWnjzs9YCUwBs9EgM77oqQR7mRpfrsbap1y
eFvIed1w+oMEyWifdWuYvASek6m+NMw4GinnGjTBTpSvid4NgG5eVMlWm2ZyBak3qXsuLGPE7z+8
sV/MjSB+7H6xABoELYcczP10rlPCk0Ac8SeI6XUhJzisyaI/TgVsfzAmFO5ohnG/h8Ia7a/Zzu7A
qgOCW0scUkKDCsInZmvdk0PZoKLR+R3ha2iv5xon9tMPrVd0HwcohsuTsY0Nmp9agNmw1Vu5yQaX
EiLMOoS27o4O/10/yuUAAWbI598XlgIgrRErEXpW6HBGvinlnGpXFaTwWPsOzljHbNP/QbOnIPLM
44/hdcU3l+bQ+GzOFBBMXcYnCgOgoN7gv82tuO/YpFc9brLb8riYibGif9MtNtgyGmh7YLQyDxYD
j1Q4AMHsJDKrmb5Qud80m6DmvcxYkmDIc53goVlPZABlswJa5wVDlzZXSDTZD1PIP8kIWqktoiQm
jUWhOolw+VIxrr9JyijmG3vrQWi9swgFwTZ3I4mdAK/CPHVYCQm6y6xwDNr+y8erL0gY3mZU4Nlx
cImYMfqtbljP95QjcpZ+MjRHKHU5bIYle0Gswq712J0EOEf0Q1kTiVhIE17sqpsGs0YvNbD91Siz
2wEiznqy2s3cyiHiJVxvcdXIhGSjRHlZm0zScwWk6W5mYG9eK7b0pemr4lN6e2UvvvAYk3MWEPfG
gc2WnaWzL5DJkLdLT/KgeOUrvod/bJAWhyZPl/J6s3t0d7dqDoF2ghKW22cKqZxJO5Obz8H2EMyD
hsUQVk4tY3oFt1O1vi61cnTImskp3o08Vyv4xPNnKp1H4F0dZO2+ZeRgfMwSK0p6YzNKbPU/OaJe
n8lLIg+scU5dgSUCoVdQRuiYTNay5Ar4cx1vx+fCGWUW+SHP0pTqGJk4Z+SheolVJx/FUefLGQeG
SG+8Uvlsai0LR+TDxEihhH4PsheplOB1inku6yLCMSuimGpfX1YCBbsiJqmml/5AAfvK9Z+9G3+K
Ag6orE5gfjG2eMYXe51P1q66qGu/2SJoxiT0vCRbCe48jp8bjUE2uchO0ciCFuN+89DebK8USzTl
bqAIltGS8Zj9pcF0MLnmMoGg9PQzYScDkIeojg6yrk6nYNO+b0aiQ6tfPZu9lsvxHNHRiYbRCebd
uvyMtV7xzlar6UGDD+nTw7ivEdpTQSNtnU0+bsOccQypoQ/QiehaL8l0bR/JKb9WyKD/J6WLEQ/A
qC3fKFyuQMdtRICqgbKg6xPrKzJQi1T5KAdqgZmy221OhsYXA9IOZokhNg0CM/eF+nKV/+peSRN/
tce/wr3SRiBpvg3e5iQzDn3+zR3kVcYSayoM1u0m4K326qoKvrwhC0LZaSeN91aecpqfM1F0muej
acM+icvq06fygOBcNLfv6Usz3Oju3BvsblvHdupqqFSXIaEQa4FbNt82jVDbh+9pRXO+P+CfJLae
DJdZBKVq3bVTmLOWo5FZY/GCgQf4f/pxHs8mVHLtfMRN0JUMKEwKbyDhokxddl4whlvqqk7YLApt
WfriTAkttZG40DA1jasRv1RwS+loSDZrXp0iRzs+pLNVhuzTEW/7CoP35Hk4NaM8kuJEMeTOcpRE
dfIHpiN+XjqJd5gj12IgDuyjajmpAs40YiipT6wGhcfHszlQVhOfuDOEbaJlMM4JxdrwwPxPzyxn
JzowTFFHIHwYg7AFgyZSUXqAWu0aYN2nnaHHP+plIXJrhDznai3wZ+FS9Qf3ffsyUJpx4GTaWMwn
rW3RAzKSxX+DCtmsdjVJpAxp913bwOTgxf8Ht0fLEKQWmhQlKCBxJRGCkBKOetOJaFTHLWaCwjFF
Y1jiIsfXzjztap8s4JTapLnrSLMukrFJwypCQK+PK5o4yk1n+9XesLykXDhyFVDJVVPJ71kWd/So
BOZI+iLfWi/zfjKgj1g5ylR8nGN328motA1tdTdEwOmESeu8jIX0amyHvzWmwEkzLyTKYH2uYllf
hpl/bPtvPCgHTFbzlasck1W0dWG0uJjfRoClHKaaQ8HDHhC9ztZxax/1pbLqkISkGsA1wOIAUESi
y3p4S1Twl+7KcI/nROpdj5xVTTdNgjo9ZOBhChoeF2GNjFsR8wtnKFZyu8r/TnfjrylhqSwsnrdq
GF+jGSW47eJB23jjY+mhzFNYtIX6r3NOXORY2dUdJ7J9ewqO2g2zv3/hQbPYraEbSGRj/cfGvFFL
Eo/t+jeDemMRvXMwHH/Ohfb4uwZxMPCWlSK1sl4sdP+/URvuOdFBxM4NjERr89dgwg3DCXj4iRiP
c3F29smAbgxu3jt7Bm46pwWMNSPC573TC5gz9OvwfyViGELzewqdY5c1yjuuKhfN9/+EaOxJerUm
jxuGkcmXggNMy4/4Pz1/V7Rqx/daJYC9UxOXDclGlAEvuuzU3yFfk1CW9OXSmKYe7v8frpncB3y4
xkvskbJeFCOkdJDYKExjBpubpd/rlNwEu5fr4udbjUyWHnP/OfeLTKM+eFrs5aLrAe+fE0BWc2Sb
4PPFrbbk28Y1dTxQ4MnYTcqDjXnApWkoum7itAZY6BqZS/8G+tAoPOnxDHW6Uo3SnQi7ojdLq0uB
Pp1g/LM1dMLSNpR41TK7pfhQ7qSn5lDKBKiaIySAzsAJ0WRe2EulHdcotAphhpwHTflFppLLARbp
pnWaEw3uJnrgy4lkyop974lOECFdAZ2aLA0+odmFF2IBrjGGJo5iwyrW45P/vDfTyEJp3YCshKX6
GVUk7ilF+ariTlhL6NEaBROKxalfGsRNByRawlgBjNJ685igVxncgGRF7QsFBdeRVNr0BClquaW7
hVQUNrgpbiSA39qC7IgUGDoUIuZTl0j+VjN32U/fQ9fATAcnPdACqmAJsb2oRZc9uRRrt9re0VTX
ppeW6E0W5GhJZ6ksqie6jklTNqWcLdTMbatuP0NvNZhSfe5sOG6ZYDF1inY5kZ1AYdE3l2umSXLc
1At+q0IT4SvWvD8Lt89Z9sUpaniN4Lp7sgz++rfd2CmegaAKJYmoAmY7hMYqksg9MLs1j8BwhAb/
OttGHiLcWbb8gOMRYEIGkKxgcckY/SHLIUbCRto2UxEt4sMqLsJDsInq2+KA2KybXjRcWUcppqDA
3fZVfsl+wKvbsueIaHZVeAx/YuzugunnD/czS2kpRPW7NkCVYhUj7OAYh5BNhpiXhRnD2e5SeiE1
UqtOBJDNrOwFeF152jb8zswhU/UIsIuRNWm6rU1roVzi5xLVYER2VKKKEaWA9s9pqN5YNNEhLVxr
xcCoHJTKhStcV71IiqtIxoaqeatQjuDOnT3BCVsdmqPK1f6y2YUnsDcx14c/eo8lM96rgYCsTpuv
bElsO62shkTCb3bAd20arVCEymuxcF7l6YAtiDBAgez7XxmxmBP6OfJZQ/AoApskFYU9pbL1HBaj
s/EHHE05piGPfBGymE+nx1NcGlHVLDi28jsMyfUi1YsdSBJIs/oLVzDGVUodaBycumddnYIUwjr1
uqfIwA3DZjmOOduSRldJFO+BpF7ylwBDorNdvGe6by9OMkQ0nU9R2fVvSaPBoKE4JjintUDiscLf
f4Hwr2FoamKinScR0zbQBLEjfVshxh+QOkqK4sbWuIsuMVFNaMPolA0eZyRBwsUmRzP3yw+Eiqer
FhJF2adofBBOvRg3/kB0WLIP4Nk8uv2H9qL/JGEhKK0YXe69wITAK29tfVLcoSGXwPpqsczZfGN5
sTVx+/p2Tp/F8m6BHWjxRM0d3u/lFNtrcTSB5NyCYAil0CTOw2DNPjgerGcskPOWr7TuB7tBxaNy
02E3iKgE6xNxKYuHSihV8EIiYK/ZoJWrLvEj+6NoUjP6N/eyRyMxoCMQls/qKwJxYx3ej+ZSVFW+
bel0qFcnysvb/l1kLkXo6sNkubB9piJGJpwjvHwK550RIK3eQy+ZO9Qye4rQOEsWa7hH3gTXcRwR
Z39Wfq4kuU4b9Yqv0nv86N8senWH6P6DDUM/1m3i+G0zdah9IVAnLqxRjsgPVwkvZ+h0V0CAHQ+r
Th44+mZd9np7GE8V8msG0MNMuY2VeEwSjsDzaMHlwsSZZKAbfWU4CsQz0z93FvmdUVRv08tb8XZp
n2QmyJHd7VeksiYY6bogK/sOh6D56Z0BjTXazyB77NPDqdnXJAPUkT5KS3fphgt/83VrcHWB4Lvp
HIOEfAVCMFkbOaKf5N4j4AjSviGSKe7Hh6e8B8O73NYuKJu07dDl/rQ6TnVkjGReWQtbFW/1V5lh
M0uANAYFyy6xLg0AEWHG6dQD7lClspjS6/Gi2F1sIoxHh2GxwwQHo7N781Ln/UEYIjaRbzJNjbdf
tQt2Swk6Y87+1e15+aysnyqBbkcWG3+QqXXYlzv3e/cvdx76lBaj9RukQKmXgACOT06AdYqjcono
aqsOeXbFgxSYl8I8h8OCqfeMk4cm94PUilrHXGC76mPOAp44b3brpKTWYY3SIkGFrfEatwqYKMvI
Ee6XCogct1GenMIMHydGZ7513IRCjd5q0h1H+hQPz8iTJzNlWm1WLqX0gqHj0OeedMWTryieP5SI
4BlG7cEQflcpsyYFsdupjnL3yAs/45tJoAzhG4jBNjA/ztonMGJ7atIdEnIlS/uw3pT8WMzeCEL7
5U/N5IiLt3bW/5epeDOMFk1tHPPjii47lfNEHyJA7ZyPxu1CKp7EfaMlNRMDQp/hQsoCZQuLWVZN
mFO3Dc6c/846oSrUZWMbE2a7BQ5RulhBnXqt6UKyP0D1mdFg4rGlPTiyxqbSZZdTlEcgwOa6rZDw
rMttFJGuxZvu0vzVuJre6MPMaQ2D2UuTeSjjW3yiGUFx4KWs5XWeOxooyybICAu4ErOILwVQ7b/k
ke0Hj0oWmHkAb4OKzObySqPi5d6q12u3EHjyPW/VxWqTToyI9VySMZ5qODqMpeQd5vElJwXGsN/T
5h8r+awv8kC3HIoeH2SRwlOflK54AotO9HpG1in+2JuIwUaV/Z87Mtvb1OTPZXXTRcIOMT58KZ1h
1I29CLASKY5/vjTKLya2TUIQCwlgCYoxnJWyqjWKtZ6WZlKvMxixn8dPzy7nPr9W3JcU7xMMSNza
2jA2UjYEJljGGX23w/enKIE+kI9qt3X8xcvKr8BQp2gupFV8qWV7gVdgahCWUsFaPxNo4ZkQrZdX
nG+ZT9hc6rGJFzJZsTtHPNDoI2JgzitaW05WcZ3A1ZQAhpeIH4bJrHpQeTPUc1N8iBDtfkDG0vUh
bhx57jr4fRaub9KtSO4pr7XP3CzpYOOvc3VuPInZ11MDGp4je6z6rHSK8fPvYUZv9bYTT2TWq7y5
N2WPXG/aM/HUfyhn/Gl3W3BQ3mwHJWV+x7ebK7Sxe2+XSSrLNh86RSMD1mccGsGqseAS+5nEnDNy
VGdrvY6DAeVDWrle6rRVKhjB5NWskXVx941owUPVcVT/Z4h0/zCJO+wKV1KMxwngnpM4qIQ7s+sq
DagUHP+ypmlBNtWtlKfukiT+RTxRNV0pq82bAdDRhhu3nE5yFIBLOJsJxY5fZzDLKEoaMccO5rmS
UboqkU3rOp+Exg+Hwc4NE74JXCk5PkS32cTXZHOiYovBWcNYmwXtckhw+mJXvsknrB2Nayl9gDw+
03j+sjNPal1PXJTTwrUci0lUIDrOFlsD/vueFzpQ+/KQnaBs7O+MWHi/PZkomlFV0f4rpO8+2Pa8
1ppSIszYpZMPkXwh0hPy7aDp3QydDgMcWVbjD9+d94cCNAtWR8D3sTcwQtxbryRupTjbFe88GZjf
IXDWd1CBV6CTcPU+jVhGyp2P3uNGPSk4rP5gT3Ky7MrJyMbSYgDWzLX1JKzV/gj7XRLgBSOCJHc6
Kew6e7Pf6SuMwdyWb0JLj1q1kSC0G6lm4+JUm5qlwJsCvFusw0unzUYQ3q7HVejDrdU6CmUTjiaA
GsFFW6daRNf+PTz0CwYwzXzOxXCZOKXCG91zpefvKy346OUnukVeq1UeVc/TNIqMdU4/6TrXPnhT
2IUa2eZKtB/r5ziQFolC0YSjQLnRZq8yrGGslxojC5uMIuNQkrUMFyHYwraTU4xbNUdscXZWaE+e
r2HHHOujRUYM8e5nzreDp0lUOilOFmmQvV1a/3CLE8tUmJbGw1CLxgpwNxjNFDqtsDD2FB5LWdB0
2vbl1xCnFTTDU3/zEE3F5eBqbeAK8HB+lRoHmdVUx2P8qI4KsDo9dNVtApYFKN6IxbHPkUxrr9/s
Bis/YKhxyYINsmljHVifTtojUwhu9ujoNrbCnbwF/cz5CjmJRxZVKvsIFL+wEGZmBuMailRxoFyD
MI75q33SWg0erEpkrXNTzOZuensFHy5gq9aaABjPF1kPiJTw9HrB4W/TBtJv/h4BkZnOqh2L6HI/
HCl6AAgDmG0CQu8PmRdx2ddFe3pTQ6+o5GkwJn+y3HGOXvyCG8HD3f2IYwz9rbCzRsyUBleWC0xu
i7JBkBQhC0fFECH9wJJ6A7Q7kf8Y7VYl2L2TmsFr6qxyY1BOgQ6Cw7Xgr6GsoE2NIKoxlosLvvuS
D7rwmLlmV4sFTNhwoXhlUpOJF+HVrWbW3yADQ/xGzLkf8qyZHcEy8qTymbJN8Ro11LEEUqZbKwDe
5LZb/v6l9RGijkLZnchpXgI1CseB/5pCbHMZFgrhfUQs5BCT5S+cvA1BNjUWh9ErblOhT9IiGs0m
yoU+pyDfs07EDtPyXO+uNUeDL5b9/f3oFTroG/d8tV6EHKdmimxMBCbHFgUMSk4EMaZbpC77bzR+
7HDbxzoXeJYjNcbLTYKZzU9kEDGxZs5BE1R7I2HgpuwXEpAMzy6HLvQattKcmZKn+PEcnHqdIkV6
L/PjPzlt7YELZ+s+i2GN4AkyPXvN9y38STaTuXnVUSDe8GrRG1YzWgm5ns/B2YuuM7QFGOTu7izR
QyR+pUe+res2aSb/RCJUMIhx8YLC2aiNUFnTElD7b94C6IGeqi+lHXr/pMv2a4befKwFNv8mmMRj
vp6HsC7UTXtW1R4nVfTHjeN2DECx9rM1nyBHPEbKn+K26jLOAV35qIlExyXl8k3w5npa0LwsI6af
TiWVOUj7ej8y+SfnKnkBQuFzIzveSBSv49WN14L+yAzAyy1rTSXU/8yOlOoLBQNTFTRpp1uchD6F
72nT6fI5NKIHmeQ1p7qnocPPYvDhAw+i2zeAzrjlqkboT5xNb7Ebm23d21ZyJ9lLKZnDnE04zyee
aSQhQsYS0r3HqVrotHpthaShfCf9NwmOp1sWXosHQxG1cU1Mj4bwXRYvDGnKu5HHqHDfMJ695kYG
wkp4IpDdxVZwJbbcH+h+7dsLt85Jeq3G2YstMMXwbLVyqmsHpoM6ciPR651lx5yGiUgBUXcUsQ8Z
j10F8N7Goi7IpQGtbbBj2Iy8f34Jmkoxa3/jc99TGuE5SVk9WzOUYrcqjwWImdtyOS9nj7Ij0BQP
8PXOsh0ASvsgZVF3AmW+LVVfNYP0XiPZWsZbueRazKFlqau2at5WxcWfizB+95bUY2BlmkeKhMOM
GOcRtus9Mid9gbDO6PLv1pHvRasLpa2EsrbYwK0SWyeaenmgSkwbCUg9cZgS65FKirSsF3ippKbt
EmPyfP/FkMPoJPM9UmJvX9j29TONd6ZhCsXLHOJA6T9q7HdD9geDhMkq0jvieWVP0GbYbTp5ED+l
g4Gab0nLt/Y/R3Prfvtzoe28nYKmnJxg6f2NlfB196OB2/NpgQgYZXuUcQo1dkEYZUE+CvF3sO+X
7WIc30oLXtSlktmYcGTlY9URfUbIFyR15sX8HRQIQyIcBKHSrnzrmP/KlFnHnsT2h15hIAixQzWz
kAaolqnaYF906CKz8qevfwHaslHrhq/thuWeXsu2KawVEpNMwFJ8eXEO/s5wwNE10G4NViifR4f9
aYt7KlVZRufvD0uSK7byCtntnSKxYD3ku2ynbMMucfOQcThhKjYAT/2E7g4hzWtrt744apA2OFjb
s0x0DMGS+iOzaHEs0cdzapiNLH8fIRNtnXu6ehBuZr+/0ONyE5qr35w8MvqKFajMs2ICBRUSz608
6vzi3ztsmv418ohJEgS+70Uxd8NEpmWkYSuVVn9eD10sso9z7HlwHVA0Qfe4DPYXXEHA1dMgAfLL
31ofak6UTaUgfVMVfl51vtKxx5EqC/9Uk1x6tovB3tMb1oK2ZL3uVkYZX7dbpinztKQ0gSKRBknB
22VNwOaNKnDcpi41g7ImMTAsg3cg6eqn9zR7fjscBsrKuMYd8aG5fWfZJi4K4MYOOLxxYhiESky+
NtXcrXxvqprhOKvCmrgnNf8qTITL8wN4wTn4b8bJmpnTfyEVsJgCZv2ZGZP99riY/YAp99uFfoh8
SU3cQJoCtXvX3OA9LCqHNUWZPXfn52tzJLSTjMdr6sK1KUvSjR1/Vb+1kHqb52I9PvFCWHg8gtl3
dyHrN/x6IehTdtoqIM4N1tpfr+DBxGnla6s5K341KQ+ZGmLXxmdlHfhjPOOQ2DI8TCyqowTw+tBv
1eOVJUuo1XmmxTW8RdqP8QUiw9q1EsqIDWzoCvyL0B3Mu49xfh42FceGxaMQnjm4wJwTFnCWI/qh
qvbsWwNyjPzDsS7V/2GzvamCWAQgarrd/AjekkN9iN+86uls5HKT5w9FpOY6PuqYzvONP1evcbqo
ejnZUf8lTSF36mC1Iyc1UdEYQSMs2irh18LExehkSKTLZ+Qf2lPw8GVivGql9LX7GcQ4eNTljLwm
OqGgmsi/PC5ITqqwMmUMlt0RXZDJL/L+ooI+uYWxBDgn2WmADRPdEo8tOfBdjRISbDj1cbTqPONS
fz1jwkkXFcEcheMDNvcFma2yIhUMXqUPQz9VV0TdsyHI7mswECTF2zV/Ur7mNFYxR9rTV0T2xoVE
pI9/cke58WJ3cIjn66+hemKL04ugiQrmv+wSf+mAGBdYhyclhifEsHHh08UqE6ExuO8iT5o8Oxow
tAjvoOerrWWWcx6S+k8B3wVZm7OvXbmeePPAj1G6Z0e8+AZz1XMe8UJyMzmOHqt4rjP9fQhZDTy4
49lDTa3JXIRNYFpUEXnofatocHU9aT0jKEB3kxx6F/WZyVXYU9+TqybXl5qeD4e02+uNHJMMG273
JygwGXxHDi8vEWypwhaFMy4/0oeQ6VCVc4oaI6Ys1oEBXHBpQNQQH09mnSgpGWwzc0LWFm3dcHQW
Xc/g2KV6Fvn1M3dKmWikSIyWbJ/naB+qPwNjXi2kiE1cZIZ36usN4UntITC6zcTregtdmZXn7Top
kcueLS67EL9Kjt++eg2vLzwuGkzuYUJdeRByKww+J5RMNvr5/bYDW/D0miWWi6DNhXiX6qHxQLLE
lhOcYahdvqAgO5fyuMtqHuMOouRiBzn4KppoAiu5sTADo0g6sXItnXPMXd2J3BplrViVwifWQgFw
qWtVFXyxRG85//KsrkTl1a5rS6Mqzfcms0HwbW710Cs7cRQV5AVRbcktSbeDLsu/enLRPfZnWADU
FEOITXc6DCJ/tjZXsk1s1DWKRhA8/nmP7dVDRxc0u3BGDOisCnaRyNHjfY7jWpvXfwS/iq/n82so
8P4gcdRsz5DZZq4x2mliZg5sY7wtXOJa74ZbcTtDEADFTKyOfrY/Wg+gooyXHQ/DxkMJDfjLbKNK
ya0yqTvVKVoVPME4WxmZJTsyhzc+xuZPQPQwfieH/+IzjBH11525ABF0LyFSa1T+t+fwvIzppmhs
ujj/fpHExfiZBWX7tH+cAnA6u05jwq/9BYSpArnXuAoErKMk+6L778I8rAkNf8HwulLRY+cmdRD9
s4geTN/tuouArCGKR0IGrCE8px99FjnHk32UIjUBsoe6ihP2hGZaUXnl+6gTrAzNDlmuemtWkQ8A
iSBUtNTxP0Osr05eP4HiSuBKQeCR86uYjE2ocCaZSgtI1bq5HlxWgwbXiEqH+9PUBcid28XBcgys
MEmvxqLVF2ECPTZX64uJmfghLYg3MSLMNcikH0Hxi+0/E0/pVpA5+eVtewqe627CcSXmE5szsJCe
jzZSSTc8cdL/hE1bicS4f7LfbpaigaQm/iCusyI/VZhNSXGNT9za4cZyhwJxpVsueLuTuQu/pS8t
geRgDGVIlfvTJ1o6U9eO3DchJcneeOW95h07exi6fnsI9q6yZkKyNGBUS9VxOPcynLwVw/Tadbym
wX09XiVlDQ5WgaLytNyGD2/CM3aJzZqlPX67MmdxizSzSFD5lKU6HBvyDqPLW2vchXXtU+1DbDf6
wDM0wPh9BRxJ04TnUw++JWFZZgb8E5zI3bkwaY4s3xDCEuNcz1DspuA2QEnANVRVu7wA6Xpwiqic
rIX6OEcXMwqqR3DismBF7GTYWMeDquBO+aRFhtXApnncMrdDwgSvGOmVD+nM4HKkzTBW0Tta987V
0rAto9ey0j4VjI1P5+N9TDLgqAzwas3feVI3QQSZESccyK5QxCcCSdx27JVSrBCnUMhk4i2PxUi+
Nv1m04+gb/rI7IM6h/lzJ422kSyOqVllDAcnalOyIR912cU9fLQsXxY8ime4L0RS49VySz44XigV
K9G5jyZ1P1s6kBX+33UIE8tBX2OdYZfN5dktMHSLzEZiLEDsrvxJqWebnU+OcI81OhBVnDfiOotV
Eys5joAI5wGmDUhAMTiCHxA5+7Vd11vamEqNt7DYyKlhPhXUvFxy8BqpK8FhHhoEo+Eu+8w5y1MZ
tOd4qweVr3yzjsvgFP9l+BRomPum3wAOymoYQtU4PULRzVnxMRkjX2+V2gtQriC1/bnGfMVRhlWP
tGkypdUQPjSLkvxoXi9AhNi8AAxnvydPmMVVlc48gsfMDhdTWPudRIGbhBBg8SGtFiRDVhDeg3J8
pMzTQ1MvNK+gF1wH4dERSiq7mQxrxheTHFseRHaTcnZJCsGS0cnFSbvbzb+cRtzTySZJuAae0TWd
KIlCFvoBbuHXU1FfhaIyCVBqKZze2O6We+rFyo1E9UCWTi8srW9gUh4FWsGCP3iam85KapeTN8v2
4bDemhvq9eF7EIUQjGIypRWNWp8t3M6lnvWgX9pLhPpcgcJCWVNdMezzeBpJavSMrBnrzlkqY3l7
1/+BmKAGibf9gYQqOEgpq0Bb2v2/L+S+bKpSUfJ+pFD2NvBMoIwbG8SHkdxMDefDYU+0UWFhx49g
SxCsB4QsDanPJGtiH+InPl9sBY/BPwQKaqj+un1L19lttfM5oePJeQuMUVwiKpXZXV7fniwl019C
lzBKZkaxHZQuCTh4xnXdAxE62ubuf5h8ZtCSWEKTD46JfpLu8c5361KX5HJP1PTqxwl7vkXQ5Fsn
BSLggio1V99CT8HCsV7vVCRAO5SoNkbt/DyrOgeNlykesNuwFUlCvhg4xg6BC/yJKpJG0xCx57AT
F7MUJ45fcvRmSm6g7jybt5iZDlmzQATdT3YJFxTxClC5Z3SGdQbHTjWYDauoQPV+EOCrzPLequa4
bPcONpylqoeegwzKbmpL3Ub2c1RfBzO/HrCV4iAg7grZv9qQFlPoLocOqNzZs3tcW21MtPD35N4x
2X7CVYGyqmYAXBMwZQHBQ0iaZjzKhd5ZTy6FrOLJndXYLUsvmEIotoJk+9HXOUCYO+zCezKoKSRe
AipxBJO0OeigOqvZfcWWoWbKhOKCn2yhag9chWbDqH1NusFbiti6SPl5h2lVqfxmgZU55Oi0mUR3
h98l9sFt0uu1svF8mFYHY3oFrFri94Ug8LYiIn52sF+R/2t6gqnKmcY8d+gytqHvY7HUrnvpcEXg
KhrQrZeImKVBacSXJGys8ev9j/IKQ84o7D+OxqepbPGFG+eAA1Wstt+aJmEg8PpQR6BWp1+4gEpv
nnMnXSYJmiyM0FG9/JQKj46FXoi+UG+VYVFhwAOlMhBnQxcKW3r98Lj1v8ZlYb3eR+6DJpsGrnTL
jnxeMZzGtDIrahnmpUZPz5WbG/OxaLDLgVdMjprxro/WOUyosmLcuyOjrsB0o5r3FgVQgyDzFb5P
o4zrMHsDPQc9QF0NL51reRgjTlQqjj11TGfCivVgMIhKOSk3AEF7Ivs09v0PpOizKbB4P/sjVpUt
RXv5OoLZcTRp8GqmRnVmIXRWePZBNGXsChAOmOCOEVxo0cPC6PA3qN4eqxE8OdlfZHrO45eQc3Cu
OM9n5PanUgTSLhOjeIbaBNoMn9QvgVJLSwaxogMrwjTaMzv+uX9D12dB/ONhVfQziE9o5FCMvm3F
11yuY7ZMmuywQcu13IVz3zrDV0pfm7hZ2avSpn0Cvpd7FKP9yrGknGs9ugyDppZ1l17ELvaNKpHJ
8UiggrblballDJczEn075OozLMXeazo78DHFaJ1aLe4Xo5kfMwSY3mS6eVElPVIOh6uOcg4KktEB
Qszmx4LMz2qzZtrd6cRuQ6vI6+KtrSPuXjvJ4OBehOaLF92aLHWLYsKqbKderB5U/yzJOYsVc0sW
6EOcJ/f12D0jAGIVgdLEpBCGoDkvW+Iw/ZHeZy9/YaaVHJ+DQXqGQY1+Y23tmBsN5QN6iT3cx2QV
DcKzLHpgAZIxoIRAFEgqOzkotiCKKPbj4uvj7UHbrFP/JSAjv+cZ1fwYMvOO+WcZ8ro7K3He81YJ
VwL4jpIQFRUUe8dzC6mfctjOkoARSqo/CepLlGnj/CTdf9LkRTkm1N+/4MAOpFKxs4QjjEEqagcE
1xIHCvNYcbeWniMffWyMeVi0fPFn3b4xkDUPdCktPEtq9PeTAOhSui3+Yqp6FpqqO4s+ECIRJvto
Pp7m4rD0tsEPJYlW9Kd4DHigaBsvyTj2kYNAV0VDEoKZUR96ePxmG3sG1ZUb1xrWJsWmmv0KiCVp
HnUBSAoV9eTnZdxahZnGYBtQXqVf2W0b2Jg1EYUgqcv2I2NSngPC1Y2U+hUORJxnQBbgfEZF5+67
HOqeO6kXS2OhM3XIr3CHsuzd+8fQ21tAa1sHH/JzHbvJ6fsVtHui5paAa7QzVtUnqlJUynK0VbGn
knr50f6YELJ7saQo9yrLi6Hh2CDwTkeqtUvJx0gmZqbkC/axb3RWiFi9M+SDKMo+89bZvGuAf5sF
gI4y1vFw6hOolyhgjh+gLd065eWJiI5ncaCVmr9/mOGO0j4o3k3DzAUzUhetFvGG9prJMLjP13+b
4IwjvWS7XUzjv8yRefKEYBQp84b0zmDDJUdTfbnMPD57HV3//GYDPifRuhL/ggvhXTs6O41qdPj2
xsqhKw/phhMH7CAIEtcYRgp8gnROurw8826kGYjhZgF7YBblhDcCbquia7TzhPmpy8tHKmCkmLab
HvX06gPrjha/i/1xszsi3jvil2qkktEsNF0vpAQ30kPFMcU2fBL8ddUa2y5EsD8236dSpds1mqtd
b78630txFXVTG+3BcpY6JVx8+L+ps55BnMWQKBw84zE/TwDO3WbcR0jya41EaxHadQM5tSa4HjwX
Pi3D7RgsZjXAEpdmCkVDEDIFeIjiF6CjXE81il3iOC2hcAN/jGyxcZM0/yRrPazrxuy2+Uqg0iz3
Iq08c0Jc+Ir10EWCHN1B+mBLwGEZoZ0vHMrke6LzfntbgJ/JoI/6heHRuJ1GJu/Uy0bKrZcBodCt
Dmb321LRoDEC1NTQU8rT4Tkvmeg/CsoXMXNr6shry8S+/shrNlFP74uGsLWeuMxdyMNkXKDWBbl7
n4yFAwagEXCCOwBj24XOm3zKyG8zQaoA43ShY6AxxMPk2vSDryvwvLD89j7AcN2Jt4LSCSSog50i
YuRI+OLzoPHvdFS1j2OpLiOnZ8L5tRKBxeaAfIHUsCa50f/bPUqdGxalJwisI8cHTgq4h6t9LeQa
OQMSHMAFEq6DukWEqqRaz6jJRQ9itd007nQBug0vW8KTcpMavj33guZEU7QQXloshTtqTJTQkIuI
nbVYPfu9rvRD8B0AEdVe+BccUDXUXTDadCt3icEd8nBXFNNZgJCGNltsts7w/CBMB/m3M3bnG7im
RArh6NPXkrEkNuezmGL92ToW2M7XYwZyu3BQpqz119n1+y/USYuu7GvmkWAepRe1uaWhDhy3W46h
scQ5/9oMkYFjyXzwsweOMgLitwomJK+IuRVxxsZjnf28OljCKdCYjb+6E6ciVocFxdEi2vMuO0i3
122Q1Wb8AljfZVOw+uHtT8E/mx+qOlgxGUHAdZsZMcaHgXReNqyj/CITJwQ868MGyKbw/mbqhB7J
kJiUUMizTu4FI6uEUD1ZZic9PMQySJsK7TyGD+2mAfj8ZCsmk4PmKraHfyknwIIteuQCpXS8tQpY
aOwkG2b/5XHnXJ/H0X014pDNkwm3QsX1uIuz8su1/a6eu3C4+H0qn9jXwVWBrDK0HVZysILCDk8O
zTrfjuvb85ExrOE6iUzAmW/vlJjdgQt+Ez5ac307n6NlIlW3mdVkwm0YjijamF5LDY2KzJNvbqRb
o/omx242ehJhQrhFEwXmCKzsGDKi/SMoRaGkO5Mb3OQ543tFPLT+PpEneHQVjR5KxlRGFI4UIIF6
xeS/sNMH/dParmwbB1iOsEVpTlYBTz7hAxjyze602S62eg5l5/Ap7ywZ5LLLJrYQ5LPXulrSm9If
eF+e7XUo92aFM/2uayr2aqIR4yuvzNSydMQhOLQzKP+9h41I0rdq4Ji8hDvAewFdEetvObpuG/6S
u9xi6TU4zxMBXLp9Szyfq5a9eZmy20Dw4Gcu+O8UA9NWHgVlUkf/Lseln8VR+n4hqVzsbxfFwymA
PPSq/VrxM8pTWKSCnmhTa23gU5JrunPlhzWWopdWe9Hll9nwp2JCNmYUEv9iNPjdM2lAwuHOXBCu
EvFqGjBx5TIMEySP2zReTwTsJE4NBCaDLAwXR4HgNRCjDJK3CFGA14Q5TpSNzC5Y06FUMbcffh4T
nvSFGDqsANt6chfEtouTbERIqHG7WBdB8jQDrCzw37stEJUOwgwFquNrxrgH2AY60o4nV7HGt0oq
4grf2L2BypFru/a7ba1Goo3ZONTJe9aAFAjQangVO+MEt8OPKKxIbyj9F8KTYnHE2Bht2gEqC1Yk
HhO6kd0wFKtocyUc3Kbrjt3+b+q+UAeugHM4UVFAz3cTEY4Am4nGaezCEqwZmNE6UNx12b+Ptjt7
w6+DJP9S3xvWkTcH2XqBB/T6l0HUDFk28Ys1iFAikJrmm9Hmf8VYMSShp8DSH8QfP9cXqmBrWjo0
u4o4rzTMpc9Exg55sGsHZDpUhXOQdJbIKpi2oMvkD7qk1makbJMRiSbrMvB+RJl/UIcOWTCYPFry
1nxa3yJUQl1EfyRe2nHABh2XuC3ZrNEzJizRSKfIGP+kllmXMa55dmKClRjuaytCbMEfkxf1fN2p
Hdwe55gUx3jqY+Q9D2JMLeiGqTj592SMM5j67tRklsHjFQn8SRpqVng/Q3paGNwS5piI9VJfH77G
OerMSnfvEEQfp9Emq8HikBjAOA94IBR82HieeldMKAIPsnT1hnHKBjjcS3R/2GaXbTcd2gj3lggK
aLlBr30HuVEpkvUE4gJHvZtJ8h6eAV2qJg4U8np2dwgi2iIdOv6ePLNACVOwzgjlNi+8fvjtz/lR
cjbEboOeoE01RycmyhRx+g4SDzg3Vph0Ib05KaU3hmT9IHXkr3p984uV/kWO2kKQiWShYNTlKgCX
EDvyADVpqtBnwxzwY2ecAuvo+G2XFhQp4AjI/cSM9Ed5nhyZeCAvUVu34Z5TUf9S7ndFn9RoexOu
IpCFXJWjmdrEFnw5ad3fumr5dmxv9UyR4qyC0wCZ897/fFObIBu4L4bUIFztVuVjn5qf8ZBboLOK
RdvwrDLLrYgOW3ZuQUURNmodzCsEHvtCUtD2W75pV7+LQ7UkpihEbj7y1Jpj8XjsNssreSTYIFn8
CpfA5T8v8wcY12My4nrspF8OktoiQqF2w0cBQ9Rcjh+w9h4hd0DmZ+mVXey/wMX0M78o4bsXVNM3
VrptBnmIDIbREzdOmhdkrFvH2TmgdU1ZSh/T/+aNvvFpabqAKcLkDNIdIdVY+j7ypHUPy3oftGjs
JdH3rRUp+NRfmGXn/yysVDXMpd5eaDh1ILVQUg0vmcUx9YAPclkh5B5oZ2KTl5hesqpxjYhgpsCv
L4RJUTf9NwAITYO2OiuN3T9Z4T0RBGPmpsxfNqta9Zt/qKdPLwvShzSLt1ktU1huc5sqrkY+f/c5
lnMkes7ITNoOv4MMcAKsh5DGfK/HP/hV6PGXq8QFFjPWV+nPzwMsFHm6YZou5Qtm9t5aGZFfiSEh
N43IKZMZpdQ0xWbVMKMXIj1oixNpRmScv4T2I29IwGsLiwzqGKwyDPuvFyA4XicBd6Sydj+yiK5P
pmyrGlJbleBLtNen3/6BL6dKJgBnB08mGHnI6SNd7tPlb3takvNkjhdFL5n87TbSa2cantFy3hFO
xzMqoOFc9onBLfYkEd30jCSbx+1fvMgKovOvBF2vnZZQTOoSzPDgdA8eCzAIZnB3RLXVMmhdrRyJ
QX9Cmn6sNDrRcjy+6QRjpTuUYtjh53ZOAYx5OFVNdE1RWPUK4mfoLnjE1KqlnNhbNXLNRqnEvRyJ
//9sFQ4rDwrP9k4+oOggauXmh9t2d1bziSs0V2DBl4xKlUiXznXTIxTDssYt41l98Thj4QnKbpQs
SFJt5JiVTPcLnJ4WG+vZSQsLwZpkQbOKEX+cNSryN80XSYndie/l1sFIxqDq2sWlPcVVGFGSYu6y
h0UG5BnOzUOgTKDSnE0H/qtGjfKU5e44odWt1fWtHUlUsk4WWRh740DnJa7MmGnYIS7cqp6drc69
xOynoCMIVwb+f6Z3hTYNSAoJA189tXEHGnOmWvMPJUqoouLn0cURZ+KbxQTIGRiJ4to1zy46oT3T
hwrZfVTPxJEC7H/L4y380Csc7IDkErudxjg31SKaIR6S6NGbLFrc3/gu0EwolhcZ0pKxptIt5oBv
4zmYTSIPww6Ci4H4P5+7scoM0mdaqXjeHzdWorOjX4/iURH9igu3Ae1/yunegoAfCtT3A1hZpGLc
xIyzwC169u/aljZlRR8sMYvFOk0Zga/2OtjDpTsxXVSEyKs6rpATd1EyMIB5ypY7VY+Zhcn7i/J8
aJor2HkYXspwszrUCZNPKpXuuIJIO5PpKu2+67pYOuoOwleW6sgpwLdUZkpQYr0aIi6QIWlRWIDu
zLJ/79vFKShwIsOsZ5rF9szncVj4WHuG0W+cppOy7C/ecCFDt8r1INAk3GDGngXzJjG+SatbHiUF
sgRU7sa5ibdjHGaqOy1u/9RXymB2A11FPfAxcfbcOyju69L4PTqNBw58hTbMyMPllTCmZbHOihBV
iaSBxmHJK9FloXEnS3u510+D2/Vq/L2Fd0QrEVCFs+lLOMXCGtounjQzWoEz2M+aiSO+0k7zWPpH
OUTegvFP/jAKNAeEbW8cgN0Icip5MEiIJtnSfSFbTPL+6CvDT27Qfqu8uufych6TU2SYTtLSs3nC
yv+nnV0OW6nN204KN1HWUtHKH2bU1eVTxvmz8mTz8A5TRu1t4Ik6ZWj4CM6jc95UNNQsgOYeUg5Y
rOeAinfNrtAu/PBUqcslStasMnf1Zqq+6m5VI4hhD95Is3R48o2iey6iKcLSGw4fZ2IMsajQztRs
TZl4EiS6Bg+cwjgnPnKNJc/MEcbY5cPqEeH1O2b0GUjbCHLJAjgqpXH+6VE3wcav2fEPAshJT56i
eCaX3wlLMHVpG6gcYWkt/IezHS3z7Ri803hGMPlDnnjaaAfwoVYOrXiTWAQrAlCEWF2HGMTZNSR7
4ZvMIoUjH922ShPv/lyDLigU5PqWgnIkWUQ1ntO7gOqmUfQHxmZ3z7UgJNUOdzZUeCsdl+DuL3og
KXpAch3yv3rMsIKUOx8RHkI+qmpwLVvZMh6HHdtg8TkeL+FKcnb83OjFSNyPWrz3AiwcJfJvYK5O
t+MIgxGisdHMgo5c+FZUAhnI0CV+ObmuDeUmSzANlKvz5VXzUG1gQnx4zIv+u+5uHEdXm6tFregT
Ejt4Gg9Goc/5wsyLFmjmFVeXWDhHTFhW+kBbLTWjPSIgqzhaHo98Sd/OpRLLIk2xwOajz2yOk87f
eLEsUZb3NPIuqiPW7qp3RFIVpKw71zzI8vU1Bi5eAYH78c7bsDytAa4OB0Qux5uvps+sAKxW+dDi
ZxEuT6mj2uX9XOY5KboIE+KmMMRGB2cpVhGS9D2OkbmzsFU4U/6O9irQJH+HC8vB0Sok407RTT8P
a9pNi/uUHgNrkgXnhyn+IkjPnaBejwigTFOinhAK+JEjNcRkpv2XCwHhc6WOWceTyOnpa2a9RSo6
uw0NRo3m8OC6V+apImYbbIHSD2J7QFRmSmJ857ctNbMOehiTqt1ov53fb8jb7gJJ7GGti71/3Xzk
qwgt3+d8wOosW9wniQg6jqoKC5e2rPpNiufgsGAjlavFBPkVG78ANe/4uINeZXVBqIbq4GFF0jAH
uJJAtisoZx9gwQx/m0Fc+Uj3dI6HLFfQi2+AdcIBR9lCS9SBw29+gd9Cm8d8HsPx1bGOYZE70JqN
wWFmH+7M5SwtXudzLfmnHsRImh49zd17wpXwt7R6pmKf5qgJNcPD+BZxkLaSyLeqICf9DhVJL6jW
D6Uv5bAigBCu9LgZ/AcsT4yzofS/BB0PT8B78y0jVTLlUZI3sIarYIVEoET6web6kfpkCzGhnEXK
B5zWcM2uPpk1P4zTlD79vzYQ/7NYuMvtJTn869UjlToAqXfzta3A1bmYL+kxV8q7vu6FWdeuNIe3
a8TKsEsLHDlP4b4AHqPddtDoCfGbkq7xTEoTvVrAyTN/bJNy1DEt+NqwaS+F7Z+ROYWL5aTJehIm
VIQxtPo2OOU4j1+UURhwPsNBadA0VfpHq8dBhg/QvYP3gQOA7gY1qtQzabFErNdmGX81g6iFX/dF
WH94Gd9tGl47guRaPlxuiq4xU3rCRhfo1J39VBydsjHyU+65hZIrvuxMLirwoxPO0OLOTAqjLNnM
vcduQKcqHx0WOkzt3Ka6TJGjLsUVp4NPXVxGK+zfwWPstIk/YbGpVh74jS8yD0c832iu9w0wkBNk
Q3jWVgAMMP8fBjpHZjRPkNO0wABj6U5shS3DUnYL6cn3wVqlxTHsaBDlFaN2qkIpSQ8ZWNYnhUkU
RaxBNZbMyNA+ZRxy0ZkLxCL2ftQYcffIYhnUv29/ArW285cS30+MGDlfV8W8IpdcNSnQ4f8JlGLu
+Ycm++0IE3nCc7bIrXhalR/iWFww47KjVmh1/2mBgCkC1GWUgZ9POzuq+KC7sDvEqrQmlXMOglip
D3BNq4SIlKflNjKtSvdUS7coIjhIdHnTnnQdKpaKPsbce1nGsyGxiaHJWSWpImjXp67DLuOfsMdY
PmH37Hl8FdcCw7MapK22X/h86DeBawBRv3+6TYVPgylL3P+z0bqvmK9H3cxyf8LCv6VTgUGoMcKe
Rt/gw/e+2woimbYW1gKsa7dKpJPP52dKX1YkG2A0LPvCVCwqNNgicng7Tbcb2YXMQ3DKrfnTkhDt
a7issMXU0+MfSZST/Ir3U+eMCEFpB1Tqz7qNdoA6+olmydn8gasehNHMkzssN2o6dVGtwbdwkvA8
xRcQcQe1DHwFslc+deXp7/nUm69r10hWvCAEb5QurODgt1p9iXW7049Zeayeay832Ck9r0OvfIPT
ceyYul6lZBSWHGoZNu7G7N+ytYqcdH6cJDVvjHWnJVawKz/qM4VLDdCEa7JVR0bPVjVDvYqih5gH
cv3t4Sp46zPJ7HeVb5QQ0vbXyZlJAW/yPqT9uue+Kyx0jbvwvpxAeC89kBbuLvotmVNOEZ1vMOPV
YTZ2xfQF8cnIbAMINtlVdZUC4JXJ7PSWQRi2pHBY9935PkujMQtuRX83D5O0KZ+Y/jmLhnaJybrX
kXV5jehq++IKMahtaDPDnA3YrFfmLjdhNhEsKnzdOdPi7qrtBgoH+XFswn+e3sUkcuaeGX7NISWV
1+XqFXzHN2BU6xXf5+u74nhNDOBtjGhvg3CseGL6KDr/nCruCMxGIj8dF/0eOty2zBVoM3Rni40s
Is5vbKBL2WAKIGXxn2Iqr07F5H5cQ1Ga3+I0shp3cxJ9vfjjd7oNjADklH23PXem1ja/AQLHa7r5
+NHat5lyhz7Yrz3gITOAu2L8OISLug/+UXRNgsbsU35ZpLBYnlt1I2sCHo7Gc2WQa6o73+2ndNBI
ZXZ9X4VInIN1zFBu9WmDsIgE1RyIPigkj6Y1YwzwCMgcWprrjWfKzMnh4rWM3/C4Rc/833QyFFrK
Kx799ReqYRU8jM7Tvjrh8jAgQEXFjtluoSc8RwAXQulPCu1hc0SxkOT3nN01rUAMuyeDT1iFeVoB
Z8R4E5CZt/FE5XV3Wh37agDwFV4TavsPUf4d1YWRGGKSKNh0QNWNvaRGCkolkGWSkv7+M4AbhfAr
PUJgPqYaJUa9uvND4HCHI8hDQtpbVyYL/OsLoVjmZfDxCWogAgx6WLXXh92d+47e3XOlY9673rCP
1vj51sfSiEGHhds2gHr/nyDibbrsgwOJfEjufAllBOhDaCY4n9SA2hQhDd3D1wOpWl6+L/VrxjpG
pLD6HJjrjsz0rBVlOT3+Zh3LZWu786XIPHHoQT8phwN2ALvEphDpWFyDmlc64p0+299N1W4neUIE
HTmCQMFUzb8zoLFCUQ5lCWV8WKai0kXEugano8KJK0lKQRE0s6wLnL7VoznNcJFAeyRMkevo8ZoM
jOHSlDu98qTjDu0Oql6xRu/DM+Ku82weL0K77bQjpHGo9YYfoyptRXOxbLIaT3zYstC47MgktA5t
I2sjM5CXIn/Te6TFynXuzGfTdkrHGeYpysLWjgV92wypsIe9GAP93HB4EJatN+tIs/YaLVvjjtj9
sjJc8iuNoCA8edanL1qwAMBcBqubmnHd+EHNNnzDN4qKyLc0RVCNy4Zu8jJRB4RatCcExbO6cHq9
au3frs5mT/HbIboBOcIa/Txaxgp4rvpJQf91nysPe8zqsPFtjthvB+MWCX0v7DNU47ld6D6z88zt
IGQs5xRS7yuVtyMmQblz0svALpZ5IjUnslK+hzp2iQtzeR1PBiiEKa0BjsraDuMsseN/XqorWKN3
kroyAJMlWlWjRPT6I44EK3JuNc4khn1GRyGURk8ajrlqKeisHO2ay+r8n/mfqIQ5vg8FGIho5ZRm
ye7D6x4o1KX85dUvGDax5PzlzcUGcJlFIgkYRwH4L1AO34DGDvz38245aJlC6/RejmVtGNigo7eH
9XUDsfOGUukGR3ahbKnHjR831supoMmy09PELXPZN93wbbPDqsJu+s44jE+uPdNYqbMpvQeJ++Mp
MwlH2BAWrzmdjqWPZa+ksm9pGFCmIVvf7xY4kQak+vzJphS5k4+OOgV/M+A4yruIQucdV0qn9JGN
LnNG3gPjXNTTcGyVlPeuHMiMZ3CFynOzyB0hK50ueOaGuPybBnXAl8EYe7hT35iNehAc9hwVuAfl
uKo9u9zboRBmRqOq+MJtF7rvt/zZBpeCsXj4xebAzoJFNXxPfeq5ZpOuZ9kUQXUVo21E8l2F2prh
dwOxoY+l2IrPvIwJUEjDA93LlihUKXdBRoquF2HzeEddJtG+vcpLZjXcsPFX0I6q9RBqSR0jiQcM
yQ0GfEYrBPOo9PKOcjpHnk+zRivK00GwBrGrcmRjV8TLuKcnMV2FmwAuJA2bZwycCRnP2G3hFs7K
xh3RZryl08e7qy/hpf22zBBxdjPBUP2X8iFI0mVzxuw1eeQnpG3EmilNoo5OQzGslOBkjS+Np+fM
8UbJoDLbbj+v9Qf94AeV7gKyCMn1iTqjlfgTSA1KPDdi0VwdIJp8GvQJAJ5Kk0Olg8Qt6ZBfExTQ
4X/rKTvrze7QSvZWTHkNB4cwkrQRdqoWkKTKVfwBA+T8dV78HSOG+VXcP89XGzd+17+92lwg7EKb
FZFbPpvY9IYP9DzmL6I3H2lmuIqx4qROCqlKyblC+osdmrvMs9Tulb7dIeSA81mdm4LAHXx7WvoA
iSEv47E5kn/ZMrNCStgTZQmzJQfZUTPRhmIsCi7JsqeIphnqGrPCi9PKlQD0tcGj/dZ/EH6Pu4O6
9uG8QZE2+5N3YRmWd2ken+jF736RREUWeviOioEYeX9ICyFgiEbpBXB7LX+lj+ThmX3W8cNOA4kz
qIiv8hvVWDBmD6SMmkwj8V31sjReaSEDmdaREq8ZReTm0mGaT3vIU5qzIUKV10GoGxhVLnQrDycm
ewdssWIY6+vCm8rx16Z1iG/vCEi/geGqWUJLXgOig3H3zyAq5KpV9XCe5FkdCKDwq7cbR2Tr2gLL
neURW4YazeP62wrnUBxxNLvPelotdYUqnjkPkfOVKmsvu6YgonFZPUyrOD2ClHmOknT9e/MsvGGR
xB0sDrN1VSrUbYjDyD5Zw4kLuWY4jcTUxozxA6yblJF0s7vgz/hHlh7vcG2rP8RKY/xEGhty5TCX
gLJbE36yzGM2Uh6Rlkdo5dFD/UcbHYyYRn3hKnKu6D1Gxm42Q8IHeC/Q/ah5Ph9QC3WmdPD1kp0R
sggcM3Ogimvv5LkbAaPzxAEMIlsrLPnX2PNeeOo5euKoMgyfhUGOlXq6gZ3XlwyP7h4GWi7GixSJ
vz+0KlOEpi394qP5ySvR8uPACEM+XoncBsthz1788P0z2KH9rsUBdyeR4v0anjTYPsiHQslJrzJ8
bTaIxDTktX1SAuIDUYCBBZs8yWbmO5frxygv85qXnrdYUxwvUZRTYBlU8wdSBIoapQ6UY0fm5VY+
H0q+KH1TuXRC7M60rWz2Fq4UlD2ib55tAGrlC728gyuk6dEiARVxkkCrcbo7AvOZwqnXIv3XdrBZ
pdly1IYUNZh1ZbGMvQE5qr4cX1Plqpwip3WoBSGB++PITNG0Xv63Y/e3XwK6BFfudL3FfAGTdnoF
YuBRjX913jKSIadBUAeWBGgcf1JuVCw+svYZGt7kCMtt9LmtmhWF9lsXAXlxfVZPUvpUQAripA9e
tQu7YiNx150SNMdNt701U5F51HibClDHcPYFwr8qyR3FyAawY0M4gWZtIuLs1potxc7grF8ptJQ2
Lz6rK05kPM8FdWBjJ9DW4ioDJmhLina78KovvZX5x4OGk14lnTn0HEhsBbtJeBuZMQ3ZGWAaGYDX
QyqUhw50wNLEOISYEeXgWSd0mYpj/2DEtIWW7wwDHqRiY90WYrRYwF4SD7IEKpc/Ab/Yu40THmas
+cI+MrkrmGEcsyhzX9sCSFyyE8zDJNzZt6bAL32LcyjYOXnJ/LXo8Bt3cjRffM2kpyQy/OK1ESH7
POWhI37Slm2uKWgLsNXy28mt1UU3dZj22cfUConK2WX9QZL+BfNmPldxLb7sgQ5j55XKrn3MGR1c
JuqNuKa+9Fknfg0m5R9WSEJ9Rl/tfA/xUxXoBAMdCxHkZDoWUp4E37Za9IFgC6SeRuxlOGSvgPOt
i/Qwqgx21bKnvPG1mXwfcS9o18y7KF4Qt7lxcliZsNQUQhyLgoDOHG1pUlNUOngvVpJMYJ3hDRjJ
YBZPc2t0iEIRCK3yWXP+/lNTa8cbMFPBswocA3pvJwNR4Pq2yDjKiAXPBeSaUGzcN5HFIT0dOVW/
HX0/ibJwUBXyaieIjjOViQgPFmvw8FEXrXzVaL74R+E1Eum331t6Wnv2gIl+Snao9veKoB7O0Vit
fJN9J9Lmli5zdEzgYQ36z9l3DhFox/K1NNfkR9t8CyRm25jJNl7F7Q5/sVVY687Tazcil5nB73Mi
9yHJo43ZfeHBz+yyy4MhSngd4h/Lu3de3StDrk3aIZTOyWko5vuW3FSXzzsa5Oh7WO9wdV4NXONI
xkUZpcCHHixA9F1bo+E8LXXnxXnMxYX88LPAw0IEwAFtb2ERobffxfIa0rUXHib+DkEN89sIbix6
MIyV0fNsnBh03Gu4SglIWoswazhW/47VdRKumsdlgLt2CdcOmqz1ulpZU66RLj31wWUYOdyEi8Ce
uy8wE9K9jTCQrLZFMtQYuY+uY9opY1QCxTf4KRvIajJaG3uUzpxPFixaButv7abqRQ995URhHn/g
LxSfAOdauGJ/WlFvFr6DtSNMyZF0ZxHCtP5vPTuLEL09dWc7p2VHI3oUICO8N9BkDdJ5yWz3XWZ/
w/edYL10taJithhIjE8XERqJdj7PR48DVtreDSTOEsE+CrRC4Z9VmM2U6HqSmWqPzhbjSDyyrd50
OK9Ppupggvhd05P+YvYMk2A1gH+6QwJu1KbAOEKwT63D5ChTGtVbLD8HVVu5kUvpqgDP0vPs1OXP
GA7NbO7m+uSG18J+RpyUHShCBCkkDJUYqJb3xM2MXseuRwhJ5QupHTWv8AdCPlI/LaWhML+cxE7i
3FbhGC2c0BfUn1FWHj8EnleJ7Y6rISYnL2JGRVrZNZz1OahI5B8cmoQgLQb8ESC+84eodrFREyrP
fNLitMLgEzEGlhfWKI9StPb78WOSIRj6+L43qRM3CoE/OyrOKeVTwD8Y9fCFEuKaBeTb5QcvCuID
gx9VBwEQF7qClRikJ5vcZp/XlzbnfhZzCGlRMdL0CnoLx3vJRdNYRIx5+VCm6WGCKu0Ewq5wWk5J
Kh9ZZ7mMp0Jx/dAs1lAnsqyWJY76IUVcnoJKzMuORtdWBpqWlq2MsKjfaONn7ua9VrW2NNnR+jD1
1qH09v8VmRTZhvdyIrbmDlOaYPrwAom7sKIrn3Zl/tKO+6iG/zEDXyxCPIyqoCaUub6Is5TG3CUP
SHYPkeb8Nvz0/Iq9p8HNRa40lPVQbkn92sgfeamPXSCK/ZcBZj1+iYgkVy9dDVAzqD0hEipSvh7x
5enXqBPb8B6V5+i/kq+k1zokLiQhI9TuqT7rV7W9ujkI4ZWLyfieWlzJFqIt6FW0QH53eSLkJ0nL
nBY4gWyp5GkipHsH2LkSEAoO8fznXHCws2FIJ0smJJOBLLkCOtZ83FB9byYhnNfsEqV2gdXo0Ir8
eG8gkqY4Nj7bAkuiqJim8Ym8x71BFCcACNO60v/TM8jMAeziXVhhXwaPxQMjShh2od37qAVTaPDE
vsnpv1/bi/vXoM9VQr/uGqtaZ8Gn1DeEl1Md0CmKPAZebEeib4q4qgiC8Io7aP9OSMvs1r+c0fs2
AyBB55Azqrd9mF/BczIPAf2MyfmQmwRaoz51HXcZhoO/MbpZFZi+M6VnCh6N99RlRcAczZIp2HXf
+YWCafuW1XeRLsuaud8PGOO5W4z5YUSnUhPY+uegPUjlUm0iaNuutcHkdhf6xgUgWw13BiuNeUqB
44zRlcK5c/xeNxkyf8TxooreEIMbeQbGyxea8Mbqo42gW9Cp8cyoRDVO4o7emtbmmK13AHk7mvlI
8qaq4oPvbvcxmN31WULU2+juCw/s5uZrsqoKVRvIyK0Rsu9wyfsNxEMy6bIH8DMboo5QgtnbZeFZ
txeiABYJxcchqxR0m+1nSLOsAONNCUjLGXfDUcIfrMGknb1nOBGvh1bEIH76sc7ov65/cJ4msGKz
2HB/X/IUgn/lkOUspXIjg8GYUUWUh28zCLtdQkUiD9Qmrc5Rx5y6xrOCQh5GyHVK73d5NMMQyRJl
zj4Sjjp0vPSBwZuaOS5WiETUh9PcWqqwJkvfXGHjrylSO9d9onYXVK65h8U43Owg4XKWj0zAYwCo
2gunJrvbefhUd7GGyFgxm8NeueHHR5DxcugNfjTCpNxjovclinop+LnzrP8LH+en9yYVWx/pWUKQ
6/t32e2lf6v+BoABcdihJtrJePqXSJ46mkRtOW8twLD//ZdoCQV6l7+VBsIXhLUxASWcsDjMdKvF
MEiSKe0v3kQT0+VlYdeOAEGwB+OSqJ+RHLXiF2Ir57/d2AJ+6F9DGSeGoeBi/QAj4fsBhdHfxXZR
spZXwxANvISr53p5elDagTc+Ep0WpZR5dakMs9PyJVH7DBTiX8aNKS3kBx+34BhTWlQDbN/WfAsr
CPl32vY4Qf+R8UXYMVgQM3hq/CLAJoa8k4vQlMaJr71DZzo5ez5brR5VIGKTbysbXWPXlqaCnhYx
Xsose/zE9bh0W9XQL/MG93i8CY6KwPyxBmG7XlASPTUG988GgHcm8WXSbipDb/+qyY4tZ2Pt0jv3
myon6HXWJi2F0UNjYyQzpPKbi+aVD5D3hdN8cN3oAuchxZH/oVzAwORRBrez5QAHXele0OeAG+Qc
3xE4BluhnHuUUEAYvoGyNEwInCQnPsDx4mwYy8yafejby2mgUYL1lXTlcG7Zy/GjC4mpPZne0Ol1
7mDnug+FeXGcxwXDIDrFO93ZTkL7wVP+eZAZe8EYkGw+JJ3YMQ3mft2qgFRN44TWHTP06OfU8YGL
Lc0acjg+SiE67uhSEIHOTV7RuxbTMrK2z0zNdn/FJ9kPKsmEGnyoanmqZ9i4bbIgeCnSDrGj2kxN
sCgqb+1XGNVkK9FTdKft6tTrNLZtzlrDiJPXJKbUEARNvajaBszlOfrZSMXMV8I9RzjhAfWDOir2
ibw65HY4NPqfjwWewRPf9oXCb9Eei6Yzlno7f5hPJxvjXoNc3zX9XMohyVnEDHLa5EbnZvmSPRCy
fzI0pZlXD1DlgcUk6CUywXfiRTwvmRELIo9nikkRglfyx0GfNZuhM5lOg+OjAH1PKsc+6rMAywaX
5+SoMeozfL8lXq2LUM2pDuBuCIOypk1ow8z1eeRwl+Jso7PcfIIbNR8ZbJ1482ZqHM6582lC8tDx
2B/ocmouVJbhuo4YfxbL9Zf2pbV0wEHlrthjQxVvtX52WIbLRYfRTUKk5gDN/5EBoD4wxMhzIT8b
KJKyd6GvmiD4OTKZTjaPVRr3kd7tl09ZuiUnLUXUSRO8oW+lNmcA2wUhSo+ZKMavAp6U/AuYfn7o
uQK8IjQv9EgMgYyGG1NmL0X6yM25UTSoJiGJuIzANxXxhLZOkuxcYtniBg3yaiM4FoURHMJ5AOf5
UZoOKigF56RTelfnGjgRZCH79ixHwI3t6qP97MvQXkbEUnaGmDOaxvLgSitVP/VzYaHKeqmifXxB
Bwx4+d3XEpEJXsDSsBcQvz7a4yTwHedORjMcJXjZU0f1C+PJhyj+agRMH3WPOlmFgY7l6U1pVs/3
TLtoUlO740hTvjIcNcSrksZvyGJv2P7L+bYW96fW5hDpnLvF5U5LR3yoydhjuWcaLKn6kqZdqmAy
hXvk+/xBfvkTpQOw7ENT3APMPVG9tJq8jaR4W9IXslqb5nJaPO2y6VCCCHIQpwmz6jU/PkwDkdYH
cVpWcHHMo7Y+12FJwaUbHlNz1OIeV4tWpp7Kwe4MRWzFahxlGTkouLcNEaSX1QwEeomTIxeSbxKE
/tb40XVyrhiru6PNU1MSoVVwGW3S0I8BMefTDpyPXQqg28wwuTzFo2EwPAGyAtBRdCYCcVjBQTCB
SnRHxg/w9vwt8KZ+2J9VzsbOyMfhDJTt2NR2QI5NqfADyy8a3iQkQ15FWR1BnQU0Y5cIhZDmR4GG
TXKuCPgIc0jmDzPtRloCEzLhUb8nK1Yj8P4bDSroIaeQ4A+3uqBI4Uf34I9PDEhdNh95Go3BRj9l
MTWAoUckJz9ZqZgkycNsI081ZIRymaI1KrusKwC/gQdRfxhqjdaGZ3ceIXiE6uCo//Qc8tj7j4lX
TPxVDhpdWmhEiu9QD3xMV1Twl/HI+al7FkUGPmPlpS0Gs69ysBqAoseXcCpfmxTYu7OqUOs7iylo
NHMwzcbt9Wo8jg3F7CkUMOLcU4Ir41RDQaLCA1OFJIq8uqeJBa3UBVINAKIRXNOuDy7FVUZ5JxLj
N3pBLUNrbzeCptF64Bo9Mb5cWkFB6aKkTWy6FN3k6bRzYw1ZZKBNk9DElwKS/ue1lugmA5E2Qjsj
wJOzwNQop/Y4mI9Zw0cfSybC0fiQzp+xsUAej+RHhJRe7FOPjsGc3zL8StsFBSlh6n/N0J47CpjM
Z616yL6zQBFddFXh5sX985pHVbqzUozCLbK3b26xAVp+7MBO/AM6KRAUHLBGznCFtMPOFU2w0XZt
A/T7GdFUqFJ9WT4sCXepnyADiHlBOTuysJs7XCInNKiinDTOYRHmX3leUXN4tFHdZS1p+eJWhjGA
JU/rBmR1yGZTZRccyNBFR84JUDWEp9/rxhffDqvIva5l91e+8umNyAyKlvoXDnIfGcfqv0+L7fR2
or5KPSknILKHUNghIsYQWNECvRFQH2g88VlYsbxyy40Vfn/hMOJ7BWxdm/DSVad+LD/HudoDs1v7
IHg0aJeFZ7FJtbk1vYQm2r9BRVP9agF4bLD7uQIdkq7fQdpXxLrDytnkrQhbvlRMKg6sXeFG05Wl
4UkaPdsFr5r2rc2LEfuRd+FfOH48aMIJS0Ln+Je5dJFSrY3iDBBuDy4KFebHiZrFnAAAa0GO/+gn
fYqQmajuUGD26K9PZb1v7/K6AD173rMVBMj0A/pIDJZlpE7tj532iQjtAYXDiIQTDMYE/b2AEhtg
2BCMt74XvgrFiYGptrpIaDbPzIJ+LQ2t+Z+tvBKaY/LudCFhbKLD3SDjsbD1rym2ejFAxI2BQTSQ
Bx4h/DOUR8e4pXmvH47avaQua89jVxFnJMoP5PB2pyNW386vDpWkxn5hYTe+67VXhYxhV7/yD00F
lBmD7/40S6s+croR+I3G9CRi1YIwtXhPSH8PtVsTbif1PV6/4LmEV99rvgle6WZVk37UsLpLsCMJ
EPqFnvugw9jBk19QkJl2Ywb99fIrccgFVcadRch1xuzEjlQFv4lKLgk2oO6ofpvKgIzoYnIjBkPa
yk4/FmlXW2ZjUm1mCDbMzfxwyOLUYGQ0wMu+H7CWD4BbH/HeytGBErcIpFMSJrvZ9GOOOxU1zxlO
ZWNS9vY7Djzp/86ILYWRZKtVjh6+tw74hTd4c3DUIjWCRh2l0qJq3wcl+c9DSt1QExSK96vWInkX
UwkghaBpOpWMpyBnCCrR4pwnzYHep+uD+US6OdEbRHWRDfKiZuwR2dUX1/wTwwXxsD8C37Mjl9Oq
UoAx5VmW9rR5loq+lhljN4OdPxZa5Zfnie476onlEBZQ2PM4GiZbn4nvSQkzlonQfxQqV3FUEy47
Hta8KGdzs1Bew8Xoi1h/6vyx7APwnSNlQjUhVb55BgzZS3U9auF3WZ1ySYOBm6IUR8ZmFcVXUSux
rl9PQWDHevdQA7ZbNGSxWru0e/2v8PQHmZJKwJ9HALi8geq95oYsD+nIy5Ylq1HJfj8eqNddKKF3
0E0e0AdvsQzQx1iW66kkqhSXeSRJ/y1zixqFsCEhgGTTf9rHCVQPnmZcll2piIfEDe3V/vdkHfBh
3E3Gt+v/TSxXG4LH6QoSNu0EMWF2eNQwVPBNKRszDLYl6yayk/IYtd68lp6Nhi1nQag6OgrbknvR
uirtUKxHEPuEKGKWKv0UKqfYYTj7KbL4Ke3ScUfzOjDR33+uTHgbe54E8NXMbmtaboj4UD+hV2A0
b6ssq1Jqt/N2a4iqL8HQQBgWL5cvk2cu3DpZce/Xj3NX4zFlL4N6JwGJ8GiLMZgzNdVcD/sgFRhg
745x+eig89DS6bTAGAyOB/vitmvCG3JcM99dColHgxAGRSrvzwM4ipENfGqls0LpJ9fc9bNYnOlq
D+fHXCspfGTZByTbWf/3f6sHRx8Io0wLweNpWoyHv0nrdgjC/0CwO4lsbDJQZslS91SvlNeHm+vO
g5Ajg6JV4BCrIVyennM50ojsJWvNykfky4ftKgNhY8bV51H9F8fcQo64ntSFJlK7r00uH63mhoey
yPbVvHz4bKD7Q07agrvz7PhMXh3TCJDNQfSX/W0BV7VwFxYFlOfIxdONSAwBj3tlgf8iVbWmLCk9
fVjipXgUrX6Fpu3TUAT80d5Ulg/P4s1b3btPV7dILmSTDMaQW78xLyCJjGnpEsdrLGA/2OsjJJOD
vrwpwinMg09cklYK44nG9xQd0eCuikV/+m6+mDvza4qIqjiJctl7MkhFCw7EWm8cyMvef9ymG0Hf
a4F2HQj56ZqbXmxdwNkQ4zSndNP046Dv5HxcE3ajptJFdvGVDUdn/WzsU88fkec8+AKAyVXb+UYm
/h8L+hpQjGGKTuzP7NL+8/AR1f1M5EIonSGW5D6n7PtaOImiGHaf/eXM6w6u6W/iUrgCMoFsGNq7
31EHJhGukrL1QAyVxY8huAe0edYetb8gIM4txVO6L7PvbisBXC0TNGzvGxeMMcx43MqZEGBHY/ze
oc2eIxd/1qLhfO08kCW3fUnF6E3eggsEp6lGu1ctFNxOcf4rYO8zKHwlQ/896LSDL3LhO3uGLoMV
PrbpPnRo7/CSmBwauYRiIoNz3RAlPIHcz7NK3RyU2kb4Wus1llwTFdHz51pP1Pazqrj4A9OkLS9Q
KqzCfvW/pHOC846P5e3Z4lQex62savg7qNDrgftA5stgIHnpfe6cbR+lBpMBbPBFWPm/jsOnsNhG
K1dLL49ufK4Py8epUCbucOvEmJXg5sG4Fs+qSKvd/cMyniIG6WdKDdeWMHKzmtj/uBxGg9fdwLta
b/GcNNdbSqiD86WkNRgT+KiZA/tu7uUbka03uc3p/DqlB2pMiU/APGGhnDgD+jVGnhSn0+6S//od
QfniqBXU0pe0FHnHiioPhATkp6jb+eOyvZB3T1l4FmjdCK9cstFaT5hhs8xtq8rBkpexJCAt0rUd
1N5/SShbWg/yjKq+LjjIgiUWlHjaPVjkNcfUlA3JkBsQUaswC8hwG+6iiiYEW4kRm8y8r5+PdauE
FoBIBB62IJIzOZXldwp07L6xlV+7Uuf1R2kV2Rz0CAYJNOW/Gt0q6GssCW0wPfzLcGXvdl0aTEWB
lkR6HL4+MvhfwYTSPMUTn7eie2RXleV5T7I54u3SNRt4NjRmipCUuqSBXROIkduDfAVRAUMmRwee
Np4C5Ck95a1tkYDTMw6GIzkgRcNJOeSL2JzbnHkB6ELVIObp6TZtb2eagEVSiLM1Hv30ozdB/Ie2
peVVYG+8EWUyZ9cKcc6yiRfsNyDqL3aGCP9kwgkEZbnzBULJjWN0c7hO6KgFK6pX4hNI5w5IKh8U
mtcXWidMrxtlzL4nVRMnKVElK/MfgDz+QUVn2kgVpvPAqDrldtGD2m7alaczez2hRQ8BhpoKLrEZ
Ce0HKknVisALZBog4YW+yRhwrpggeYXo0i8H6UbmZR8ptqwzbIC+egN9YwpTNKfdr3KxpVNT2C62
u6hNLcOcQnFKA8dtYPeHE90I217uXgl3wJRMMQvX4Ha4fka/24eurREp4Yf39klEiBHrBzILmGIu
9fhNuhskAl8u0HJ2dNkigtLSIWm71joPoK5eib1cc9PUPkKKImabaM22AWgV9KaG9NKZ1NK79yeJ
5bTXayjpLX0VcmayQQOsepZtbT9mAnGEs+pRzcnoPKDMayreSvt4RrwvR8FuG08Wyvd4VaA+ygMs
bPAeuTCmbLIwpL8B7WoSUEYqr5SKltBSKEWVDfYWMg5KA2ZXV5Ggv5E4Xr4xnJBwwlJU8nVaEq1t
9GYXxor+aAJnaNkYk7aXBv7VFCywMpTK4jEaVfRAXqUAYYpc+Q4AIGmgJpGrVPXHzcC4V6gCkgD1
WVT01Y+TL6Tu1hlNk4ta7Y7YyWiQJFMbfciXSRgrnvikX3UJyV18FQFmd6jza+tHuM8ng+KQNMr4
+t42VBpzg5LQGddX2ehLteXfffyGXZK+kZ/rZogkAnsmv78mNJdgk+3gS5HhVw+iL5y4cm/rH3LR
Scj3QFXiFKZ9xXyop10dXehweWojAVcetrcdi6dmVAY3Npzvau3I0ejoFDyWD9Yaa1BK54yCDtep
gibtvyCI218/QmgxNsq2r040k+7DfpojSUomvDmccEJIoGzRD0dxEWe1Ev69ArnD06s6GJM8IXeX
m0STULbSsfSWb2HWyBVcNMNHPq06mqPwX4usBDKcMMdt/IE+qsiptDN0JqkmRfG77ZFCiys3haSS
nctyX2DtDLR+T2kc6fRABqY6vy+lM0Ct1jBVZ4cXh40E2sHurZyuXIUHY/KZ/TSxiF3eFkt4aFK2
uUcHaPmyTpvEv4CTeyek3RAZp1DLhzN0HLL1FcfZHwwh40f8fgHG0deULpfV+vluNIqpSlArHPrU
wY3N13Zt9RcWRAt3oaKuEZK35QvtBXk+bpnAD8i5WLSTpcGqrZV+7fFu1e4s2zwOPq/zaD/2+RJy
SlK0chA15pMIpDkMeUZRTRw1U9V74BowcwrusGHyMsiO/hx42URV/d908wRW0EXHKEOVvtzwXPqm
iIashmZjNgpyRp7kbWemSdldbj3hDW4S/gY3zPFSUzgSOArN4UiDl2/UyV928Pc0YzhWq+aMwKPw
LojvYnfiXNqKHwYoRW6qqrazfWu717tKjzUSf88MKS1rJCX2hO6j/vRwc9Xp6pky6+YBsX+CL06S
TKen4NruTVNdwiEn4IgAmruvkRxkVm0wBQT1oO4+3G2UiJOy1u1VugMeutCFR7UiC6/qiQEC4BiO
XWi6dPDVe9KaHnxKmp/Zo9aGmCduVuaSTiE/2HA346ZGwUJgUI5VmU+4iT0S37ScGj/MJVguAAI3
rSW+o/tVx1S4K6lZ5VKxGmPtIAerfktEz7MdecwzMIVraqtgFWrO/F6haovbhT6GsoYb3muxc04L
EcxtTDrYU26ettII+d12je3xRW92HQOpbIhGfT+3qKV+lrneWC2vAREIf3yAEAfPrvNuFaR5uj+2
KEPuof9r0hjl5MTmAb3EuVCGMiBzxFPtqaWKZFb/poh3behxSdsZ3V1QNvNNI9Swn6xplgu2t/eU
wN0XLEpRSM9/+05f0k7Y6c5JlvfIc27u91eNVmGrdl3JwCSmQMLxgFcIfclj43v+utB7AfG+Di3m
3VTUeOETvMWIC7XJJObwgWac91W8kLrGKP5k6SxkdF5NoRGC5+zZviGIh1IO4S6OcdU4UfQ5Uwi0
zPjmO/dm7LD3KTLzZ+SxIJ+oh3z6H5bSrWkpi/SffSVwqzfob5KVmJ+CLMakbMQddeUL+s09aPY/
mXhD90MNuvSH4kQX8OsF+aa7QBOV7fDPhr99LwXV7HupZEU7O5+Udq7Ye7bnz3WZsAzcHjN5/zYp
OlpbEwHye1NPmz38uC9UVWpz6yOYCcuAEPTuWuPo39E/09RHb67F2hemxKGIdKFsmZXRetIxV9re
0Hb/UFvJSwyk1D3L9Yz33WKzU+FFxoNH3MhnUikXg3ETWwf6ePNv+/8i6VQ22ZdUAqOwq/oH1Dkw
jg7m3xQpmP2NPuQyk9l64sH2uWAdkkd1uWB76e0i/zjeSzPqJAvMe5W57AtLzaU8tDl2Tm02Fg+d
xCJN1sgSOzjxBqRbtxOrHhq0zn0lh6KL+BIqQY1H9nY24HpmdEyaZFbSFEJoIX7b3rX0RpzSy421
ycvpXHy4FB++yRyrthJRsG9EX68IlNDlTbIPh5AqcaYPZd8Cuv8EBVrMxdFB6O1KYqQoaS110+IX
/i/i49AvRRNyxyGTE7nrlbL6RLC2fFiG/Vz2YyupE6FtDXWSo4g0y/p36C5A2jRRSy/D14kLinPt
fypam7K5qJSP6b9UuH81kAj+E8GzaSRs8o2IuvNYSTmn94N8oXhjo6YaqGXcGBMwelfZRGsTNH2k
kyWHMQURXDFpBTmIBMYkA1vXYq/FK+vDD9zsSepV7uDibljvHO0n5HRCEkOInyJGb/W9aO5mXDEO
muLK7ATsDPIu+RnGyrgHN8eQBZU4k77GCvjp80Iofx/qltllBZDAjFwa8bjUZnp8H9C4A7UF3KQz
N5h+SGRZbSr+BRU9h9oCGWrbDayI/b+P8xD+hMjceo9exwfQtfYGNmcCNZpdvtQZ8P3/TMVTuNWp
u1tKKZ4qdO99IwVbd4fQjdnuRsMR29ERngFvEAy6mWmTFQIMCXtnnaAdgawO/5jG9xhycoAGeQq/
rsWj1DD6lllGuopQFQVJUPOw4iRv3fPbN4KojdIz+aD2rntyQF1k9QsxtstHlkFnetC5ZU7ZwPyA
XFN57jqRerfgo1ELmZ1HAfnKxFJtKV/c+H2/dREWKX+Ws6JzigPYM3LBrV/cw0QaSZZO1q/MZZH5
f/+mjdBXV64PcA+NKfhTpmf90CE+g1a+E3g/U2OLkMexNBJ9y4AXRdBbZs35qGwIjN57cEQhjv4Z
LV7L+6aTQd3EmHXtw+KGGQgf7SDhW7tab3mZCtJNmC8VovcaXR1rfRBp4f3u03KaUBFQAtauIOMO
pGyG2wdoZ1ovzVT2OHlJLE31giox36OUW6icxyYAdqN6p+QsCWNlhkKWvYYMDirOMUCcoe6R3THL
GucZTp56+/qP6euRzvJdhp3hJeaUSI+jQ9fnqS4u/J0AIZQ8eOl2hDUDmxyMcRat81AVybcZ+Qdb
Lk86bAdzZq23L1VGZbYtC7ziv0DszaGhzjLXeku57LgGWjHFFsoiT9xuVlFdB/rT9+gwBzsAJHCK
ACLM30+kh4Dl1C71cCHbuhWyBAHDJlojrzF9fqZKaMQbqIKe08dAvjojL3k+rD3bMg3O5rJkY22k
PD1uKq2y9zJEcCyLZebKNGAlWIaWiHA5n7BUc0XygZXtMlzt/CE1w8/dBAOOCiyyQ6fAgVORqWji
jmq7rY0wL8ay0f9BgZiqBQ1bf+dW7BduwoMBpQUg14tOIuheh3nGkKinjiNW5qr3bnZKl65deqDh
wkksIMMaN1HQLdnCbLqVb1z6ws3QPypoOtCkeEFQb/UI1IWGCe5mDGqX0wOelAfkuHKg9wUKEimH
YzJoA+wuU5vEICCMwlCCMXgl4tncAlamh2x5p4hT0FaAJysw171kgy+M9Af3LzM04r/ZAfe05Upj
q7ROOvNEo8tu8/mKZT+pYTHMFqQpMjnGk0UN/g+amMSi4LGMePwGGFStqOzeWses2mHqHFagQCHm
FRiaEgP1iss3imZwnITQ22GXRTDiCaiOVp5NZ1JTJwTDXVl6IjN4zfXw9B/bxXV+2WN5rhD5WMTn
WH7T+YMctfnPFh6GkJ2aXu5ARGu4EvLQoWMportzWrEFNFZOE7U88o+qNLQFtmI+Fb2cBHMVhJpR
WDXe+ByxLq4UEfZxwvaGoJNzLEuZxMsyIB8IAmhrLApt3hpg0jikA/E89TC4MLTpoKGuEo1eFyee
QATMeOK1XVZKlFXpObcwqDQoStpP+2gX5klTPENUTJgSo4VPHqFe53UoxmdkjPBXw/MZbZW0gxTA
vVOjikKbSPaeO7OPIy/bPB8u8rUpDfpgvr8mc1gmZlDSm6i7vwQXLFQDhxuMEYAXqRcYg0HvuSTP
zaMQeHu7Wb5TyYmqpMRcf+ioNHz+ya1TX/i1S2CZObI6EVc1FFy7l6/8qhRvQWoOusLKVzOTBy7T
hmQVFW9QAAmJizTDCFl7wCaSakOE/pX/GI8Q42bnaL1CE9hoKQ2N5B7Lwpr2Z9LsE1wg1IT5Fc1I
qJ4dV/bOG4oMn49RIVTU7O5L4fdz9u97qLaC5mNsNQLyMwqyubjxhQMrXHca9GTEwcnIuSaNgrTs
fga4aQYthIHkxZYqZ98TuXirOO4rV4K54wirIq8Yvh3i7A+bm8bfaPaqXa1qrSFGaMmXN4x1vlpc
CO29NV5hNzfAPWHjkij81pCgUsw+RRCKaDLDH4AsKkQbGi+lLSdbL9afL4e/0jw36zYOUJ0iBUNK
V3xowI965B/kEZZpuZk2VcsEMbk/0pJAXq5o1VcA9c7CZ6CIb99GIMCh5PJRsPer6YZr5RAD5Bzc
FQrQl+AlkIGcsE+WKybbQGWMBXqOOtx8RGIMFCttwfuer7VIlyQXVUg/dOxy1pyKKwVSfHj94DOK
WcJHF9qFCxn7aGgY+vf7jwT6aogTwWTGqU29hXfGSjXNDtOe9ASl/11VveUs2IB1/LnSOMlr68QZ
GjD7ZJu1xIhH9lL6pilj5cbDg4oOrCskLR5oTJ7agqZG6e8PpOKK3Ak8Hrns8dX9iqGEWOpdeCJD
jwIxb+GNs4vkTgbPrs325gq8e2x1dK4I23Ea2Lo1/dx/8homkaZeXA58g2yGaaD9VLXo1qFoQVr8
GVFlWwiVtuF55p/ge8IKSx/UFAAHRGolkLcjpKqKIWfELFruIDPas6nRrH6AtjmTvRzY7o5kCwEx
brx9d2A05xygI01/7fJ3UOiEymDDkzPLy4eQNZs5eMB2pPTDDUNPTUbb+vt9ZSvuUBstRrM3F0qE
mJFDW0gRQyAmGba3W8/peCkavB05k973PrRGRQbsra5QWNU2wjZ/6mQcF2XLJKirzrAbEtNhT7lI
4oDhg9A+rSRUMmHG0bbEy6OWZcpL1mNBXLLF+PvIN1TRHzn3mfh97Wf5OO4CBiOmTVG94R359w5u
JGp7Rx0Bu+Im6cgwVnKeIYpA1aO3uz14HX+lH8/4NR/ZwkPrxXjPN9MBIG4y2+uVByrZJ+P+nRoD
64AHU1zJuYtaY1pYR/1I1IPwfXVkZQ467+ap4X8Um+NwgX1D/yucycivlnFDiVfpNK4kOZ8eFHhU
NoW3EVgVPg/0dKnolAAZbbnT/PK/NWSRLcQEY00Xzkx63e5QphuOmAnq+IEnmKPsQsJi3v8k3Zxw
CJnb88MlzM6BRr19kWT+4yj2UocSluBuTcDHYNGCBYpvnfOq/tyKW5/MTY7E/uiIT7+YrO3MTX51
HPLk6YfxCM9gK+30xZyZubOOQD/qfXhRi7fzmlv5N3m9wZsUP0CAimOcmFyOPFJharV62+4WrjWH
Dlg/D4Odinb8cynEGm9s4fJCKV7X6sbcMeiEAWUvdsYnGegGovCj75rAKGumgw4Y8AjfS/dVMAap
K2apwMlVp1uxdV03nv6CujQvXJ7sJovTlYsW5i6Wub6J0Oh3ZhuwELiv20FnNqW6dcP6VcB34tFU
2NZkfCHKwFMyJ5XRKHwOlqCLGLFqBiXG2ADJXQWBd/ZHx/vlAPYrtcRooemAkQrcVBUL7FrU0aly
1OPGfLu/VWjniTRQWLUL4a+iUju0iwdqghQ6DL3sqAXl/v4B2rnW5TjybRImWQ7XQ92wY+pOTdao
+C10Mnkczm5bQIBYDADIMgpYJLuppTaLrOD8VwLOlIMey7ShDfF0VRf6zsNZMJ6iv60KJuNHnSEr
rn9+x/1oPYEoSoJb4bc73i7l9nt/KT6MUsiYXT8clQQxT6t3z8XfMLVz3WpfZH6l9V2IDjD1zywM
ottdFnjrI+Vp+lGErPrgMmw/J0SmMs2yaPc7ooMuHcXshMPrc2H+dC0Wd9aYjbxwiu2l/qUM4T5T
VX683Ro5+RY5s7ECTJ0okdWjrTMRVKLFc3GoxAfmR7XldQtpDk3agxAdBPcT5VaHJ6mgIPSnmO83
50ErPmwTiGK8TXZJuVdKATLS4j5XMbpHKUtYn6grG6wX6Jb9swpo4kbPmOgPeVbrZpaC9LyawP4A
Io66ewzHGYAOKQqiVCdu5VaE4jXMzKvAestqq3FB3rJw0cBuMx5K5rnNDzgWr4WhI8/eEVKlX296
jsh4JBAiktiHPXnDka1ExuCXFCzNr8N4Bhae6snPzPJM/0AmDqaRqT1lzVUJ8lUa+ExAVuyMUY6T
1Gb7kbxOiqFCJ4KMwO9C4ISLZ31icEFtYhQ59ErDlgCvE4P2jTbJH4iLf2YfRolHHt03DBbfGW46
LWHYW29nVwZQjqVTYU7+oAkn/xPvqtCgk02G9NGGfdQN6mPcKSWvA+xl0MQbJAKhC4ZTAQYOy+C2
HqSzxqg5iLOiIHxSAv0fiCAjJ4QZBoBzTmZwECjAN6ELlrExVV6fAR/jYTuqPaQMbTixT6zUpx9M
b4M6oGVFdY+x4COCNpiQRVS02TlGWzjChPi4K9GP89hurO2zuuQoH9uHVDTUXhJC48EzaXWQD3vH
z1MfFI/iHAQ8jJ+fdZK4jqQmTH1DR4e36MoyGu6kVvzx04Qt6pi3flhq+R8bnYeIbEox/ap6NfiH
DKddtLBG7WSdFrVW3/4LeI3lr08TC29+3CTg9k03hTxlm5QLSx0srucIh+WvEJ/TipCzxwzty6OA
eZiRJ9dNZDSEJ1VH2PfJ9t58SS7NPGFAcFc0sqROpH2OS9657DwYNAGQ0sbY2xxKZGGwenvDVFgP
5ScVEeAiHeDyk6lNHzEA/5pGUNEk5BEs12WWQJr/7hm2DuQyNxCd5wXX9mFdE5l7bxc+Z7uaif+K
i7EJgFHViUEfMNrkbh04jarmYMl7mZF2/xfagEP22tEzhtbmq3ak2s6NN4SVNAnurOMClBSIX9YQ
fDsLnAlwY6GoTS2cIjfeIXWitveU5rSVIDOtT1LjY4isUBSYEuwB/hCCgzGG7eZCgLkcM92p6xjG
AVDARubgjY1rGZ83Fh1zKPaqLs59BZB1erf+ERAQjA95xh+e++N24ajDykejE9TyKkzb631zMp46
THCULlF8j6XidasLZ5wLxWKvF7Qcl2PmA3KWs4DNW1gIdreBg1i+wqMWcbbNLW5feyfP+b4UVW+m
qjLhdaasNpAKupb38pAZNyhLK9SJdVSji2KHtrKAob4sfOltoSOykiE0k+2kPmaSvTP6Cne0UVZQ
633519ynhVr4FmvJ2qT+YmUjqso1CXcOyNBuTI8u6efcuybjG7tDF9P/9ikGN5iqAEBpPazSHeC1
rcotj9R415edGvjr7MvSdUlnYPFk02U9Egxxl9SPLfRLE1/31mcVP2DeF0L0LdKH9jVjk2fy+5z0
YmiYRqiy2rd2AJh874gTk6QiWdsAkBsTISoIz78lLCS36AuDr6m5+37hvBigYElRLYm6gZX+RdJ8
PKbvuXOuETzQYUUck3FGwggpgpUA49YtkY05Qj6X71JKJYpkbYy9/3pVhfeuobIzy3tx91aGXGn0
2e7CXjLWUi578HhoWRB/cl7EzxyDu36xXLSt/6eQ7zRiaJ7jOPiA1HxZ3XooSwl98ZW5JxF2PDFC
NZkpIup1RzbVeH+TkfpAg5FnUq17WMytceqoj75DdGw5hjugSzwk7Iqk8RcwfRPrewaPHIoG99I5
hcZRjy6uhJjdKnLJQ5sdeKxiyYO65hcA3/5n3yunI7fIaFICggWbqJHtzS4Dmc+NlIuT7OweJfpq
hy1hRxgVIqiZCCDOkqwaWBDZLFjl1LzokdCU5JDFjCvWSmwijLIT6/rEwNA2kK7o/NgWUSZx/2YF
uOVtryBQgZsDFxSFsd3QisaI9byFFJGKT3Wy0TnGwo6biAXlE0Dw+PE/BlSrGDAWL1BNZCbtfRez
r5G2a8cUcO/cQBWpRpEXvYYiDizkDFgNKRwDQqrApsXg+YcH/iFPG4y8OafuqWcOsDsn/AOo+Bau
i7YaPDs4u81U5pM0/6gEVpFCXx6Esu2hwlxku3Qn5aSZnmHEIWwrKZUvEsPGoFRneSUm00tF4M4o
RDiIOQWyzPgMlnP/YduNZjoALu28sN4x7yAqoeInW9gx+L87hGAyDzHGjgCNgI9eXLefQo2FmY3d
51gY8m2ATav+YH5ef2YNUxoAhoO18mKEtRBNh6/WpxV2A7bRlgzYmhlIdNet+cy2Gkb0W66/Ywq7
IMYDUvUzM0hZYb/NXDmmDyEw+pRvP0y73WEzs9FszFuOCUqcneCdDta473OmHqmb96HVZDvZZpx6
h16uUVROPHFFqKuTTPgco4K5yuoZz/cexbVo0q01Va4THTrBlY8Z2GUqTpqgSzbEWvwT/kLgnIF1
rB5U/orfP9hmh0kpKK8s/4g9GHpy1hNrwblr91llp++HtjOdI6N1LIGc2nN26pPHeOOjMKfemZJH
4JkaF6kevovQTPH3viHoB+4MC1k8Rn4v6njCuBW0mAsHc44bifel7B0CFyv3fp6nsHOZQIZd6sId
yzMrKIcxNHSZ4bZ810mCKKh3R8bzmOutEnLbuaeYkMN6rejJIW9acT/ClRdKUu6fKtt+Y90+sJBQ
7NUeClRCH89M9iyPuDSmQxADs/p9d4qx0WGy16RUEPUs3442lJGwiOz68Wg0dyUZxyQS4FIIIuX/
1rG6+2IqfoOCOqfEZRKXvSqixbivR16JOSPcmK/yeCFM0eDGXUkY54nswhFE47o3jAngyn14iU+c
Np1+nKMhOtEMqJdgUUykbeNwXOAptE8mo34OpNTOVeUSmduXp6ZBFaAxuJz+Dxd06sHAvBMdOALs
HcD48vy7YwSEKOo0Zp4sHapvyxRv7Bycp9ZXF+m2dNQpXUStM5uciOK0IF+tTWrBmnLTNs87E9pl
1F9CKsX5t4QB2xYbrDAAjTnXz9mzpGYIsKH4Hz+dD3FhHpNEjTMFUQVGntg9msv1eUC9Plu94q3p
WoWaMNq3VQGHFgzpksorxR8nOk57Z42XBPh8flN+tg6pu2BVy1jnpR4avK1Zr/X5Ip+UOPl+b60B
J+VZ3ECmvMSEQ6xLJagnkidMORV85TAm/pksmCIsjDlAkMLuQfGYg+3YoKKedxqiMCKC5/2GZHe9
AxRIB72YAA+5iRbxRknKA5bEjhAKf7iNY8BgqvtAdfeR/c/rG3UcymspfH6advWl2jYIgBmU3+fS
GZAb0VTOtW8RxuQan9iq2W6W/mzwL9zdANkvmcq6+cuGFpY3Rcz/VbZ9VnszcE0wjktAWwMgB32s
wWkda9j0u2mmM0NL3XaJAh7CnPKEVPBilFDwBfnGO1ftTvthXilKzUbGPh8WUV3Ltscux9tms5Qg
OqBj/o8M8IoTIVrHchvWpEYuDn66cbjilbbCtz05E9OYC4BPjMr8DN55xoUayM/xLCdTS46InPRA
scZkMCVlbv5jlx79ZmNkf3vjeQxR3/Hxe6M1fj/8VyoNwQf41Q4Phdcn4obQ2II7aGC4Rv+mwR0/
sCuoIXU3wVvmITjh52xlUonE2j2qhHFz1EDY4yfLHm3w7j3jRdjuvhnLQ8R3JStLF/VVBRPSUOiW
CsVky2dzDueg1zdFMDqsOBOFyLy3Lkr5itRvXDETJUsnrpGrFyWbMIX5kKuLUVKGHfnjNBjrLZc6
bz3bTffp+LL87RVlxtkMyK9Oz/2egIBQhXP36JmYwGIyIbaRCf1L4w/2SqadSrdkuv8ODqPmX1yj
LKEgIpSfdqSbesUx82TY1/nef3l+ymdbNvCqu/z6AlXEQOr5jqze5QQe/VUnPnSWu/iK/zzHB9bA
NC2Igder03hjOy0k46m4QZeNzfwkQ14Lo1wS8canA0YNQd7FkUdOEkS75y51AjdsvvEm1DBxZf1Z
K9HptnEqKADkiuehe0ssg+Hs2BEiN7ATGM9Ymz62RVvY5uYJWVTvNuGphgDaBjAP/RWPT2NeJWad
12xEg40HGAZVvFblv8xup/wSL2xTzICMnPfxbuU+RfZSRR+ZXTwt7e+oH2n18zfvdNjs6hFJq6+N
VO8tjGvPhBObYgsQuTPrbHvKYEqW0YLdzpPI/w0XTC11On5eQsM+3O2FLmQLDh/tOq9DXC+nIh3i
Qk/so/GHCMI1o32JaxsC32Z4YZ6x8Db7DIvCo2AudmXYap4mWN4DGUkk+iKGBGFphX80nw84AacD
bZXyPD0H7DtrLTa/pOJBlDdop14Fcmr1eIeBGor9ELotd53N4Etx0ED5s37T08oNJmWd6rCxPk+q
g58Hd1UPel2VoZYheV1SGW6r7lKdixDAFkRCLH1Kup3shG9GtrbuQtf8ZGSDzODo5pC9LO+arwNk
D+zOH01+t71OMQLL485N1nRGl29GMYqqyzdR7eBEMwAf6b2NCGz8/RBYuRIHfSGZYWuXQPynlH1F
4JTvhf1xyAWG1HjJ+xiuABfkxdi0hdkFK6YsQZmFHr3HASCYozGRsUyBPd8D+aOw0rDb2yDeqI05
sgJB2D2pciYTTMHwV/3lf3wZh4rNVIrPO9eUcIIlFRgy2eX7mC8WjK6Gpp31TdUMGl352PLrDimu
r0amG68CDS+poMRqKH/GXijB8AaQpwyQiZHo6DqiMbKtePqEY7iORby2wgAwq89kdAtmqcBUf3bb
I2eir6E4vx5z4VRBzYX7yQwb8K+Mh3Pwa3YUlppHCZ/0ttsWfujv2awxyR8SgkO0MczKexHvWClG
GhiaAGmDpR0qn1qN7Cry/9IBZfljvuNBBsoUZhauhrxkAB0VwsGfOha+I9SimsZCJN4GY0lZ6WNi
DhZ3iQ/T45Xi6HbQuWcuqZSHMS1pZ58tUhMIeCvnNyGWTX444e2Du7ZKQ+wKwaRNhrqlVPxvWRxH
0esJF1wbWQsYOGyrOX+WNKZU7DGdw+kBLAvH+17LmY73QPmzTE/qlNdLOPO5PTWdfXeq/5s2mzQ4
z/7Ux15Z0rxsi3tVkwOZYuZpbRzipr3Q022f4ujl6Fd2yRdrMp9U0TCER+AfVkrvUXfTRZ3Da3g/
e2KhuZrUNhlQsQA7FZ/cptN61Ek3FlCko6alfxX8E0vRFjoGHzA+VWx4GdiN28QFDucXxHh1fwS6
lYai6Fhe3DfKAzBhPDXXBt676i71nToQPRO9dw952pN/eJ7bom+WEESHtYWhkqUy3nbST8p+3ylH
LJODs4XuwMJFE5AiLKEWu/L6dCz6DKo/1nzwMNywD+CM/J+ULkg0UuhkZg/C3TaWyYtTe82LJ6im
USM6+SLvi+52JcM6HYgJ+s4bEKCkTe2NNBtH9XuTgvqGgfrTMpXtOrK14UD0oxu7h6S0GGglzhgR
G7JOE0SEBFeKB6lZM/QzH/YjtOlxtcW8RtxuOClJE7p+3uCoULMdm6Hi1puNPVtbpYUAufcgVbK8
Gkt+ivz90urEdi4jjQXOlCZGx157afWxf24Ub57GqnoYpeUz9rA3Le641S2dpf6IFq3c8x0H72fs
h32t9IZgI0CwTLRvR8HgRUx081UpZrKyr+pRBTFwvr0SEaCHvKvDNoaOMzU4iRukPcitjCcnO3Yv
SoxVdMA68MUSSVsifK4ibduet363PFg1svSPf3JUM5o1xQ996UlFj0iOeX/HiYGmucEzwAjgPuGe
AyWETKsooD2f2YciFImtzdPdpAXRr6Og/nIZW+6+9YgmbctsfZMmALQSj/bbhfK3zQNJVm7D/GRZ
dy1O+gaZJIsurVqCrlZDX9i2wwvABjzkz8XMq6lfkaQ4P5nPAbBk3Mw3d27/ZKslyWup3zOxRxP4
dDbtEBPGaURBQ4Xa2MihqtR2x8zyaokj7NI2lCIJlExH9NsSSXLUzZggdiSfScoYyPysWsKhRReL
9qnmgPFGSyR06JDR2MKi11ZbT1uOzXMGCaQLXQFutO44q28XOFZm+JR66qV0Q/bAGHpGlVBj5OBX
ySxWetknhbW/ptl0sKx5rXB12ga/kFp9McOtaM4jbTNdYqOuqv5m+sTGBFI2PzV2uxHokd19h29k
LizAP9XahXJJvyhnKLB3ulrMm4XSvV9wXzK9wCMfqUv0o1Kl9hzppFXrm3Cv4+wpXLiOLadOm9wm
txwZ4n5J9cB1l7zjJKxBYp0rWO91FqP3+QsBxNDd8y5k+rii4vJ7JEczxfNPjP818a4yb2mbdVR+
KGpUsB+03pGa52w42xbuT8/8ySzYMDmNNHeV1CWD3etwwMbQvVpkxG8EnlmDGWkQnJgB4aYw5ypq
o7Ow1MpaRZmN5TnWrKKNkrVNYqE8qMfAi8UlZiJ5RQ29dfCPZbNFdpBjj7XKTQKQ37zfgRQDBDYx
Sz6JCjJTFLwqezAEup0bf0AkwVi2a94+ti0sG05uFR3YV4L0YpOJILUCRZUAo8wlmcXpSi36Oe69
qcXHKsTuCQp/eMeCq03wNZK1GKRyfXoukHYVIlv5Ay5AnUR2fnqpbCQqCMRBFhm+pvC+CjrjB5aw
IZTbXn73+aQ9zyTqoMBgHg3MWcRQr5qua13COAekb5vZf+oQglbwnqSLn2xhez/abnpePRQrpKH7
r28dXBo76NAgeR9wZhCqYOUQ0h3utrUnlZKMKmAtz+kaSFLxoLaqzYitURDhNIet8pjwNd3e1xsr
YIBQ3HFgr/Yuiero1E6PSh5IpDT4Hmj+luRFhUB7HQKfkuHJUaUBNqg1u4zb2ucPVZ14h4EpbNOC
G//ebGdRRcCqYF7jBRy4XjN1N5tZh2mjCwl0vOYv350JfZZrCIhxPe5K+bbZdX1qxlUQqMzWdvMr
CiWkJWHOsfMh9b9kE3uv1fXwmnstwwdgm+YwQ5UpFIKkoJvciWASUZrLXUaloDkKXAMB3OxVBq9L
EktyNoFQMZ0ZFNdYAaBFzZEoQjvLlRvxJlarYPrl56yGP0sBoPkJvONIxMzpywO8CAjGP0NodVIW
Ahdync0h3um8a//Kx1qg+ecFtjACBDb4QIkXIADm2K2MSpwNpcVMVazL1VMeVpcQake91VvSbU1Q
c6xLPHHAGYZ7MErtI/5dHheC1/3aJJ7LJrYe4DUATYDZ9amSeQa/Rk/kCvHxErJowHWgbgtFTyMp
5YmCwDexr/7QsjOEdCWV3E2TabterQdrlw7jqK6N9gtGaFttbzPCi5KN/qnT9IXdrligI3uBlHj5
6iSwdpDh2wus9hgwJY9jAzkHM9UvPqwjNBhKx6JvRtche0ENS/Z+VwcUL9tJK6n+Yd1b0CB9gmSg
0kowNadAOZ4Qfwh4FpePCi+ANadEpou3IiVE8Z+IwU+1qnngRXqKc3lMsDfVqz6QqnugFR98v37k
xtQv/C4XID0D1cfM9JEkf76jf7k3pU0lE0N0nwAFICWmrkNDt71LnPhC9rc7t4SA0UgaWokTfwkb
KZP7SjoQrNlEyqSawIcGIYiLMpEzJ//t4k1v97L8kUrFbMFYkPS6ctZvEDgpVPDKn/nOyUnIeUi0
BIccgAhMRBmThcQDefnk3lnpG8Wx4Wm355jMPv+LpMJwZfjyWqIGUn356t86G7sF0LnVmDWNSy6T
yc908W/o9NJUapV0lqGGUYjGaRfvtixf+lAzyyOdK4Wgu+t/swf8WOHu+4KZppWvmUh+Kc9Nvy+g
ujgk87x0pUypZFsMMQCs6esEj5D6FR4PLzAGFu73Vj/pgwfudlwzQM5Is2IVPDzhfeXXvfoQ+9dH
q8vx7PQgaHwh3xKTUiW27iqiEfmQRFP3I1LwTBIkXLiJ0aHGMK6Yd+yb5h08aARunMXLFxLpDJPd
/8ZZI9vGQrHdGNWA8glOKuC0iybqnTP0+PWSR0WQRmrlFMMVu85HM4B58SYpOfw6pfB2q4wf/Puc
PiBMTjNCgu70Ht4wCdTbm3u2oDOq/xip205p7a9ClanGjbl8lQct2YhpGQ62UC++8FQcZxUbKlG/
ae+JClRHc46VFDsVeBfYv/WaNlA2N2nyd2UkrXYm+Q/wHdoD2ifboTkyHEiymiz7AT/S6yMCHBbb
cwnaPkcP9YnrI0kMjH9W1gVLI+1J7s/WDrtapbJ2VW0Ssbrz+vCSRuTE+12vbDniHkiWOJly6nQ5
Px/d0a9kTpifJE1JIZLjCOrHN05zOsy8xemh7QmsA//k4khBNCFGZwTeDkXbkVJqHD2zVUZJEHZB
PhPVyZElxCuky9WdaieVwDsRpM/DILaUtReP+y/3h6XNICQoi9fjN5986AbBb6KUIGo4ikhJh4XG
AZpCt+HJAxgdwd2XZatV2h8DuiARiyEE7fwh4iG5HITtSL7MznuuVhYs6ik/wxbNMiHI0AcLM3I3
9oFvwB8Wt7GOCI/64tVJUyl+7Q1ytUrhjVxBez1XYP1jbax5ONQ/dnzxC2OLfLFejGof/XtcnLXn
9UB70T2wNdSMJr0tNXxqYzFwvHYIRdACbKwPwQfZLJI+MF22pLqpQyDSBWCae/7tkog1qJzGk0gD
v/7Iv+KsfU35UysvDCv2NEYiqa3Za7HqvQ9puKIIS0C3jFmvKWEka9dKRuZ/hk/Epu/aQkDpyA4j
SnLZOYO343iXPPKBRByxMvD9lWcAg8os0wE96Ekw6Hld4sLIynZLZbtyQfZgvDnLU6SZcRKf51A3
p16fzBOKVqR9ibSVMG7gStDgHOrWvco1KiDPEfcxLlu/MTnWvBGrQK9i9oilyT6CnOtWKJZUWI6a
MHIQL3xUGX9+OLhDOzYCX8kC7F+1XiZWT8LgValBye90wWEiW5d62uV5luHH+3fM43+p+aBRT7Pe
ghhN+ipkZTjr7S85OHb5Qbktz6Bwp2RCyQraH9EruBmeZ8dSXuLgAspTb3HO+zSstAuwZS9T1uxE
Q8dLl+V7pWxRb9BNCavh0sdcWYYtiydDtLaVLLIZQJvHNcJL2w3lmHGgL+Z3bmF7xujJr+u37m/0
uDiUpKGuA4kllcZeOlKBlTnI1bc01yy0dMf4O5J4x4LsllRQ2aOe0ylSLWlYdVvj60QKoNHx1Gga
0OCdL04usXEJGRvxloa1DLTJaBmxF57i+ZgQ2CXMD3lA8I9c05BocsLXI8O+CXIzbi6rCvUMhF5z
4i7c3MevFEQVKcq20T+jCYetUQngqAzTZ3cpPudm130UwEK8Bq3VcEdhW+eWFfr/9mGtSdeBszuY
0TP0IQe+X4bHEmUkDRM/l+VdAPgrSpSPWaxDA03hAADStpyXCMiH3JpXxUU0eZTWj4Zd9l0aVFSp
yuOOfPpIlmQKkT2I+BzIwmM7THrsT42JLVSK8iqBp+nw7N3UGpPG/WjJsp3QXLZcu1C6dBY0KFVj
waycdgCshBQaCbu7hqN+YseS3mDylb5mrzlDlyM2D+Z5h8afC7A6XmQF/iZ0O811T4+OosQT/gMM
+d6ZMcEjjdE4bCt4iKkM+4id6+zWdTz4xbR8xw4yaDA20tWmyQT9/Fz8eEaEuCZdjEfgsVbzxKpg
HkiBFP51UpmEqstODmcc7gyjAkaC6Sq+805z7HSsGRXhcz+6CAoMyg+DpD3EiU2yjhHwefjo4McT
JBRL9I3PWXdfb1bVZnDcnwGg5gzdk33R+JSrAWF3KacYV9EpGd7UTUaXsbPgpvWNEAgvKFaMWMe3
g4b4Pd9pgqhIyaLaCG5NpcbunPWdMFNU8XCDK8irH62uM+SmlQHbVAdwPJmNo3i41DXT0VeW70ty
Yy6jTwHqoWX8aWWr2mMLbEvg58abVsQ9bVRh+zftnP3BAZQWQnvAKntYaYfwU4HNNNCkmzWZL1Gq
ghGsjOvrLEdk+/frZ7G7lRI1Hiw5wUSyoA96ptuSHkJRJ55MNB8mvIKZaIDk7e3e4AozM2x3GeXK
352CgAQj95I20uRkRJo4GRZH76ruht5HWgKOW1tn7i4QjCMZE5SPK2uf1iyePw7QRNraKvE1BJKO
qF+RLOHp3SslbHcPfrv/v81rk2BgwkPR4WIv3IVKLClfbwpV4W9d+jRZouAMyacCUcXzXp4K686c
PuBC/a0BHOxgyTG1dAchrfyJNbKjnPhc41rT1z+V3qtIwYh40Z/dPsXhGIlC0zsz5fXEhNtdXVQU
icR2TwpOC1FYQl0lWEpldnrHKro5dI0dtQRVPDdMQvHwoKw7uAv5txMdbfrfecScgN7ny1dep/z9
U23v3MH8Ofwzp0nEgUhORJTrtmo5r3kSKy6xTbBuYobDqCwrKi3vowcrsobdOD6wincHnsQQsZSk
motNzOqYszjgUu7T614oO0PNjHCSuWVqZrlRGoHdwt+BVFcq+nUn70cKm54o3ma1Fwl5mgkULCUJ
/nYLVvYxRPzFp3TmbYzVywXUn79aXxyy5OcylXdOpLZPwTW+B+sDavXap38RwpHDuuOLgrWj+qxs
DteJFYxo2ehJbff9ATOHR7JDMrifo4GEV3i4xHP+c8lA9B+ZOkS7L2hKJ7yzkd9RFAFP9KYbuwn5
c/vNer4BPeI9h18AVDGw+F4J01eX3XCLWPk7XLlIZPdt6tzWh/P3+diFBRuvgYDyWLTxQl5LlrQl
bPYGgiUtOpB3WMcR76G+imFYNwfEED/uWg5vvHhIPODbnlVRuJvp/zJETTTo3ST6Kkz3Er4xWalR
gV2jYAA2NLSeqGPw6hOhHh/s7kgtDI6lMEeTOJohfrdSdG5E1iQ9MwYdIpnA0v03chnHaR6fzxEl
ylI9iHCvR+t9kmLVrfp2FYxClaCMbqqHg4r4WEvQtWFifpZA5rCpJoxWxjoB2b8uMxd4Ke/fWJwX
RrV+l0ihl96cON1q7irp8+tlJvzVpWA9tqBrIfqy0aliMQdXTIzJidJF/Kt7w19Z9kmdDIwMR0wb
R3+6SXKKUmjh9U/EsUg8QCwcEL6VWI4eIhgYYROpwtmr4rMqvJJXteoRortt6ANSeWyvk5wy3Gj+
FIsi6/fkc7Z7yMNjleFNsCD1QkHRk3GLu5qVBCjmJ3hJsJQzi+TPvigIkKAt8b8Jga7BfTlKBMAJ
gcBv3DH+wUgfHNclwSQFXFKtu9H9o4bcFgO8a3x/CGmDVL5qkMJ63l4ZhqY6nu16X6NdjyCjEPua
Su4kMLBFGDbepdqWOGuIE98LVGSdAKMJavqjDfegzVFJFUFd/STQMX7blMed30K0SobSV0Fr3U94
4ftRiZhfPWha7MINeNdZow3UDRJ6DZTvb2vMliP0xaFp38P9ZvQV0plDAKQc17c8GPHNlCNL/nYk
UTL0qKyk4fs397c2y5knrUJTbV5NS0zCyQ1SaVLr75Dne+yRWxNNB3Rc4okVAoh8WNvTtU71yOVn
sv0DLsEA5UwbYsBXMzCqYjZjvy+Az+mXvXILP53p9o1T1M1JkmkCq+oHNIS7f/LKIXHj4rxzsLvi
gNZxtNv8DMn55YRC1VoVJB7twtr+dmLZ3aCkiSSoK0XutG753aUThIozJUwyLP+5mbKWzC68xcfe
1lqJGv1ea6vo8/ngGMKGy558k6x5JimZOXQAIOWMGR8g8aAE7GrVvn90EmFtyBCyII69xsNkmMMU
mOWH9cuhdHw02yHww+3vjOWsu3yAQLUrUnCXua10fdXgcnv6G/DGq4iRc8THwcEjWueljkTNg04f
CfGpWv18+ISmmXqjAlsqLAHDB47f79amNpLirp/6YIzB79TIlO7/pizo5q8kbtL5679JfrhvF7mu
VeEAgyS1rbrLDnKLzY2dlRxn8JldqFmb6C21Oc6izLa75rq7Tx/9d2JxrjNVIR8GBsgW9uYuqPfu
4TgDwePAzi7c7gl3qtf9j/7WE1Cci8US3cLd0QTgpLw3uwqipG/N7vBL0B6fa8jQyWDIHwZyiyuE
Bt8hD6hyIBMEqZ83AlZRlmLDo7DZOI4adv7ISWtkUdx7ZArL0TU6h60utuFBAnL2d8BrEzV/SBow
ag2l4azTVOj2WfAsLH9o/QE7vYGZD5VimLfQZbHGW6QHGTDhKixlutqh/dHFiJbrpCxUTGF70aqw
wMVPuElFUcAeFYe3GrTh0SdOg+6DNs5ad55tTkqtjsO+pdLnoxTQOP7jVHemX5CyPvwwNU32ubaO
tgqt+HaBXZEY+VNHFRXYBwfYSvtiYFNR/mP2EEy8kKKJFmwgYqbMhfY1/N3X9b2QSQ6wTWgOT3Kv
SS+O016Z0HX4oiJsj0n7PbHlWkT7tpNrw4BTH9Smrlr+44Syaf0tOGDBKjOoCLRFuIvUIy5KXqY/
7hf9PUvRaG2/DZmJ7jLLJjsd6Uj1qyIxLhzaQFH1nAnQyvEcnkGts3hDH5mTdLRPop5qabh6p5HN
h3/JM5+LXcg7nrO9rVyNbI3hiN58v7Vnn0GcqMzwzvezOrdzZS1ekd7yDdaqPjdniNEzly/owJtv
94LStpggvO9XD/6BdVkrrDJSFwtx6055yvbmeHC2BbwZCnjz/vu+1KPg0BgRtK+kVzHtJ/BliLLS
qTuNOqGPqzaXFZ/+WckB2baZI8ZppFtF2LWLxJKiMTQ7Q/Zq+PiKM3SjGszVKrhWiE5DHQubvUwN
1L/Q6nO01xSAuIW9ZVUTWCIUe4BmW/EecFIeR+P48zf7UtT8LW/wPgNi4nUWrFZR79R4JjByitaU
9M/ilC9ZW3Hu38/ru6+h/POxiSUf+cvxjhxT1RrG/tp4ToA41J7rQDbPZJ7jJWvEM9rD+shyY4S2
KYbjVW8EPCvyKXHeQw6LLXLWWERqT8GpzIEi++zSgkNF29AbK1sDRm8/13lyN2/7D6oLu3Gw7UGH
pNSsxOqD46xywnlZuPlwiWpJAE/JW0d1c96bEQF5cuJTEYBO8omcoh5unXCNT/ZViSvG7zkeTCyw
55+yvfSEzfpclUtWAfF5XhQ6Uxq5zUsOAH+cTLrmKhRYQf0ugVHrP4lmWRnToPVqCSi5GwRbOoMK
divYdbQA+nkmB/QAGtYn1RjV86XmpOpVnM9vQoTJzeb8kIeGocnabGKKJqj9xvynX7LKZXDlm7j2
YoyMrmk4yzijQ8hlOAq9ONzrggyjoI5LKEtqJ47v04t1XgfaBUzDjWfOCxJ+xwMAsStWxvZh0uJo
temT7CpAYu7naDmcVk2WoSHuh7cU0PTXksQTFwkBf7ObhgzzYYgeWBpaXOKXqUQjj1ZMBZc05d2v
nLlXMkhi1da1r+sK5bC63APlBH/dB+q3BymV8MgDBQu/fH7dkA/xiJ7AAw8F9VQ25w8eTgPrb4B9
4ZqStx1rg3HBpXKnEgKUs+CyqAn+B2/LFuA7em45ZCgnKM/+BSGsYt+9bDKZbnndNq3SvARGV3ny
Zg4n22Xr8Ape1hw5ByT4a8UpqkuLgwNLCYjawtFQ8SFlXr4XIQgzZq8BBcEsnDcWZdqD82D+Sspb
nn+LgKdNT68Ni2gUWl73+U8oB8uRDgGcI+ydcFlfiXFVnm43XZjxjOWy3G4S/d4nPrWYgAwOJXiT
icb12R4E1cq16XJb3p8cXDiuG+69EeEFhjQXE2ckDjjYcyOEC0QxG5YDgrpR7c8J0P6DkYtnpM7p
2O2ZXAmAlhlhzUJnO+SrD8+/ReGTaM8/Hcp/5T8THi5TYXsxgkYVCIrQ8+P7KRgucrCsBI8Bwhj+
GfZwo2Svq2jB0845KFyS9+IT38liEaiDqpbt7RKZiAQJYAij0Wj/vdvtCA/W/uK+bxnNDjtHdeI8
4mt2yW552wgp1a92TIan+nD21/3XEedJG43cd6I82qkAzLaL62lBQfW+rFgmUpH6df7Hi905K8Mw
tqAMypDGYogiOQSlitqQ45q4VOmR3NveWG574pDAjP/Yh21GgrINL6docNMD8eQV63HDh7ZHuy1E
GT5hXjH2k+mSDc8n2eTBUpe3ApghLIdVIesFnbs7lo44g+LS86XGnTFZo/qWy6Dzsxs3WCVPFERA
ZgFDZ05dPuNn6GxytoSaYML8/yc4cuoG5EeRv79J7z/9yXTP/G091fA9jxvWX6Q4NL575xXbVs4j
Bm7GAdZnEUUOutXK404h7vr4wzZEzNKfR+Lzw2vw9X/zfjRMciAtPlKzB33GFLA9jrcYor9UysFl
5cHw6iZ21kqG6FjkooTZQqp6MGMbpmVfMRHTl6mmrw2hOM6pye/nM/g/+28Wu4buuwFTIXmr11Cp
FQqIVuaXLMOBsNSjAqBMgMh8PuoY5KlqMx1NuTEx1VIaxJPi8M2RjKKArUiXFlxhc0G3EGy4+Lbm
8WQnBROzmUM0FRdaNnAT1SlFznpdXvKEyQ/Jgbrjfsg5oJH2+nAhNVR0tyKwm21wx7V+JtZGrMlQ
i9RDhKJvkYUqcA/nXXid6CcnCuTC6zErFXM1LHluOtBMCPCJLU9Blg+CrY1L6GJ8T+tEgvkc5Gu/
VydezrezbmN4AmXXwJOmKSfiXdxt02GIb52MBu7wmhL8M3ZjHTOEKZvWYIfxlUJIJUzQ4LZtx7Vn
EOSBc4A6CejbujuIv+Zr45/2SsvmxZ2Ga+fegyuUrwHjC9UKxzZBcKlGPJX3Tx6GXrfzMip5wSKq
rcDoiKHyHJ4t+KOSU1LyJVzSlsxeCpOXB1sWeHuLFaMYPqwT/UYfo2qzH27QQ+ED2krctLTjyDtU
qSI377fTArmpjjofToSYY/UUftP3oBhkUCmOO922swrQQRtr6SPv7yvVVl30ckby1o/effXppMxh
xQ4l4b9VgGpVjtyPyJdXBotem7hOKWuQ2cIYWY1xZ/ejl/viWAe93ysfVgOqQezzrRslWse2Gda9
PVls7qlFzU86RtaHMpUBhdAIKbSRiQAtgskydFxzzDzuTKn/De/r6KFt3mM2Lm7lRoFgytWPMA1X
71opvXBNEOJu51aay4qwtLlaU0EYY9AVCeXTvqxmOqTShTgNXdLJvUiO/HzoRFJO1juRpER9+fsE
VDc0JEdcBMM1wnJ7KuERTZNc93UPu+Au7wy0Y5xFzg5Mg7kaKo4XnX7T2F4dDDf6I3sc1EG7Ri0J
VnewA0c/GKDsR8jKJN2CtRvk1E0gCl/mwMNxtmI5iTy5Ac/g3KjtMwrqzKlpkanVPxk9nDvXSfeB
CrcmgFICUmJNoLVn2NikF5rjj21Vl2DfR8T7mehcxR9IFJ5oELORSOfskxnM8Gbfo+KC+5vilQk8
w1ipkOcJHo10qweF/1YXfd3zfB0ntD9/1FO7nMpFAZN+hOAJhFmqEVtAXzHnMKWfp4ysUP1MEauO
yvxzSCg+hUBejnyxQfIhVSyz1zn176jMrGwbuT1DFm8ZFR99BxuSR3CzVDhdKWi9UK53MHI7oPrV
p6bx+juzYJCrNEodAf4i4VNyyoSLIJBvpub8WGuIPVz+OWe4OBYaybiH5ZOpeOsTqCQC6GAnxEY0
heIX3F2yQWpjYmxSKfJwGP4zZ5893PlJzeQ4k6sjglnyXfLoFXLJiDqWyCbrxsw9uF9ZIRbICW2I
XCBEyuuMfbnNJs7xC04hHjozes2I6wRgk1StJMfCrc5sPnwQutp9PiVoaMQrZHxej4EXHKyhzzUf
VIBYubFfecxsR7Z5/ndmuk/5xqSt2nhA5uocXd//4WojODK0iNtz3KqOsRfu/UcnAqC4F6gNNbzV
+t6W69DZbQwrhuhfXWz6VwZsoDFGA2+dRybtvPpVuqZkE4f7UO3j1Gxr6dFN7FgiMrLeRtHj1Tse
M6SqeuF0TIIwDLbbcgK9bTg9rciGUUN+jp8tSEyYJqI6sfuYy3NMsRZWOxY8rr+BFARIHzS1Eadv
L6q5FmkIPZ9VaHwYMU3HPaI+JdyoJvgjh1n7YpxXqjVOVrUWCimoC5a7D63Q49vn60uFE9aF2CQ1
KenGjYnQuXcjbDWTMzLvm1j7PogJ3wzua374obQh4YcRBSQH369hSbfPPENArAYE18LOZsKz7pyr
Pf15P6L16SAszsqPfLeHjcV15JJ9c8QUcGJv1YiHTneYCGjR3PBUbalnySAuWTAXuCJxymF2q1c0
QpFLaqpmlFC1SDzBeDFUS4OvE+0YM1eLX8fUB1L29lYy/sh50Q6bxJ325ES03V/sYC/DRcDHL9X7
JlT+AfoBwdL/XDaKTSVkBAq4AkX/s9xnExW8JGXhxxwvfgjTMzPLyRotNfdig28IIGeNSYi7AnNK
7VODNI8NXT2Vtr/+L4YLtkyXid3iZDru01GW9BC3roAhjzBz6tQYGnAcv0zAbWqlfxcazowPBzQo
Y8eJPYzF6a4CaLzjG3y9Aj9g2daclZWwVDsg0CE94Rt2Oll1K+gCct9BEhuBR4nrNnvh8th6r9ib
Z2E5nQWHHfvVI1UXPtAErn+t4ybfTJZYZn5+YfpXpqRWt6/RjtVDInBLwnOQ0ywoqLfiI5v6d/W/
hNJZusak7RNvlPJNcmdGZ5J1YWX93Og+lGmnPzOcsyW725Ihe+FrRQpdLhXOtH8ROzm8L0YefGqO
DdpupG4a02bQxiuJicPwvupjbHIRVYcgKAo8V6h882S05TaqtvY2yxzSZGIcrSZ4Xp0oKKSeYRD2
MsuvFufvO07J/YYknqzMVFSujnDx1nZqmGxVKYLE6HjPQmAjuwd2k6AdlAW1dIvvp6SQdolkq9vK
DdZWJEufPEcXkhfXNTlako//WShUyr7tY8sDzFNr6kHkx+4xvzvmiouJdBQlgX1dq4jBC67Sv0FL
qvBGY55ClA8BYGb8+y6RGYTb+3R4/Ymivs3c3EYsOZDH+7fU7VkKMUOnTW+ClbH3wFCqoX4KEzal
st+zRfl1g58QxyteISsedf78c/9yyE1TcycNPYrX3AfW6eMWFnfBboDJswmCAZZOJ+ZE0/edYrEy
2gfnn+WB9UgBZIw6ttemFrfKLpBW0QEle5XRsf61GOllYvxLm6PUA89Uuv7n2RgDLNlZ+jKYN7Wj
13cXktUbMlCrNZUFPcJ57ZcvsxJN1Td/au30FfWkjSMLlP/TsDuKc/czXu03FbPOfGEwyWrw+mRO
IkDNIzyBnhutXBGB8zBP/gcW2oQ/4x+rP06/n7PqIrizWGVPyjvR/xgrslPqTxXdLltjCO6q/twD
+bxic1+DQ/tUDhP4HzQSXIMeA2Yj/jGZsaFr72dXJHPdvK9rnyv3PFj3ndHWU/fkpOeKaDRVBWli
+GD2ptNACVeQnECl/MDoCAQ+S8AJwlDm9DumKvLD5gkTUsa8U7g9BoZ818VHfXcgdKJed0QPRhed
1v6Uqs2KxkMzXt/3bGFx7bz3llgJcidoMoINADEJbVf7hPWUbfxlvb/vdgZE1fpNKwrxCKll5A0o
I6dTwhTJTpH+ALwZrG3g5QHKzC3dXaMfaDJjppRXM7d7lFlR9R5Lp1jK6/Ms35e+fv3gT8gTLLrJ
Sg585AD4H/V7Xj6NGYUjJ4Jenz39yMreEkNuM1b4fcco7rgVuhWSMxLXUd24u/B4X1qA6TSflS3d
EghPm9jEmaI5gYPcX1TVhHwmwZis3xglazGxtIk+pqNFz3T26PDzMX9jnW4O8PN8BlV8UKUxk85Z
cQLR6ekUBpfWECJ35WqrWU100FMoQa95FOmA8tNqPjYjWevbPY+ZqzgNpgA/NTPd3WwrZDMhHdyF
CH/uqzHYcgkqc80Q6FkHOtlGnmdq84kg7yB9SJs3BlBBw6cyrt7l2A+KryOXj1f4EsIb6IkItYU3
bCaGW5pPgt10iZT0LLxO3FCdb+gBDPYk7vyhRKFsCnQVGp6H7p1EjHGMh5e/cLg2C6wGmEp99Q5K
NsSWVi+q3dtUEz5mi1MqUMw4FQoHgxLKsvFm45aMinBQQhqC3UPYiSQ6rZlON4lUf2x5psZIrH+I
2rZaV1AaANfmZpItmCmykmdVao3IBMUFoQkGcPWw8E2+yoOAHTIwZ6BlmMxjURoyAAVif0mHSF/J
SFI7ebq1aJNPyZI7EVs3x5/iHKflLu5pbML0pqCGwmC0cdb2SpncXVd1JNlt1maW4I8UYB/2K2GL
Gi8F7aHCKiuyC1V/b8hFQnDBdfgX4Vq+kIAnNH1EY8tJzhKVmO7EKyo2O0r9IMOE9bxAULfuMnED
jVLt49f8zjMdEnRfZds3GHMxfLR3muE/lzLRKvvSQUZRwtNMxo+t9E0biBVuef1akGY3FL4GCY9B
NOfBrRGNjPnLIIiFy/IkY0nl1jskyUvV6NbSU1SVBMeV3f4SOWj1f13wnMg7RmRKFaBM6Je3XLTo
3/iLNLuBK8a2z9LR0juN+fivuCRjjkXg28Pm4CMIaY93Bu1BBoGKwj9p+efZJRJklhyHs0WAJoln
1JiZGrVuCKdizDB8v02foysAEAs7g3DyV+nqmGMqElGn3/zBQSVrBZz2ZekO5m2NHA4qT2HNxP8l
769XCb6Qu2hPsoRWcFOhnpc95p/Gudx1sc6qN+m98jhjv++hHhC7D2GO8VtmlnRwsvlbRk26MIqP
p9irXOwwuz/TZ07QqiX1lOFD6scp1RgpmOosW+n00Jm7y6wJPHa+LekaVQo2Zv9M7l49wy0NP0mc
qXQl9bUp+atBbmuVKGCm60PUhtMJldT0LdQH/KOu54FHvx8E4spknmi6mt7JIXDSfSRlBINFr9Oz
MYpaCmSiOqVyNqUjci6h6J44ym8P4e+EeunanoXco0oBFjBH3xjXYie5Kyb8WUrY3VqCaqarqWYG
Jq7Sw855HA3J7RrnSKitEZwpO87BEpXxzknINskG6l/4NeJtgi10akGw2Y4eD4UEg5w2J59vgiB5
875BEBBILM8Z8p29X54Es6m2DFawm1auxKDLzJ/H/XXYNiCRqdhR2YFEk57pLJgaxBdyrUbTkBJU
JUxKO83R2S8rtJjNhhKYqotfO9kY4TnCVq7u0TvYQQGCJQ0fA+iCfgt3MXljqzX5XS8v7G1IAzeA
faG/fODhHxv8m1BAY8mSbS2wxoKEbSAB4dE7O82bhNoMrYICyu0lXDidRxzaxheeznb/LFyTCJY3
o1xBCvtfP8jRqzNao+SSxy0g1lC78/qTwGIdPxNEDOTVLvYxn/6plBPLZt+l3MvgVh5QOL+FRHDn
BF2Y29r6bvgEFD1HHw2ZMlfD9CsXTnNJNOojaTiN/ArmW5iudZ9bgLrt0gcdbQ/ql8B+orgsw6qd
Pu5qfj/ppQoayPX+SUrdUqDFc+QJdyL3BvlEn8qxYS5JtyEmDOP1MeuTs0OVezuD+xde4fCQdCVn
/KFu2JB4EWcefuACR9Fpf7PUQXAHyo65RdMGFSu9k4l+Ue0pIEgZuPJI64wKbcI0BrmigG/lwlAP
O5X3MvWqcvvJDKm30mVZX1DPHG3xL19MbmBkwIdWA/5FBKTFHttDwsopm513EOF0SPwjwJPwjDOW
O3e0iHU0gY+je2VPPNh/aKowr1OfNoOgzFmO/I2llpmI7k9b9E2m3wJhoVxHpQpFVtjGBgYw5Lq8
7P8pgB6tVvZRDEu67CzChtFgQNJeTV5WKF796fuIZ4/Y0Kl8UbAFIPJ1a6Z6tsmV6WOqHwy20KfY
SkbGK37A8JIZ3ZakOjWkMKGK+6S5bbXtQ3IRWUzjmywxAVsuJ3EuFCRDvs+rbdpROPpk+7WXDwNz
y6icTG7VF0hu7gAlJKe2PSsTyVsQubXthIyREmEEXJTvEl2L7ZOLoZruwU8Tlp25DoY+Qlq1Doqp
9mFf910Vd5eoNmcQgeFbo21h91qpluo9axvbtRmfqYb6lvit77PBv3jd+Z1uqKpB7z2IQSXYKx74
KjTq+PAPA/46b1UN4/73EO+Q5E2DxvJzA6NT4s+w3pMhxDmmWV1o67w+95i+B6rvuH8yTuwv1ptb
BGgY51+o4yc5ERZ3GKrlYEft48g0qhT7jhN/LqMlOFol7Hpyo9rGsNSH97BSHbW2Opd80mq1ILpD
XKM0LijprF5vXHDc6bGwLCEAX55LLJm00F+poUlosDGe5QxapR/ma2tckbGZfFP+XP72LqnPEyYD
f1vubPQoBLixWokiEylb5jx7qeo1iJkjKE8QOoYkl7bCxMfhBgkFfTdL5ESB/e9QCYMCVFFGGwAO
JG9Xpn7iaSc6YHfQiDDe4YWsYZOZ6pU6iXzBAbVwaLjqwKZbk2w6MPEZHhv3mo4AyrjCXbiHhu4b
cQL71rkWgGrHFcMhgG6Oz3H5/z2m0ccM6WmLt9nrrdbw/LxUyzE+jvsMJeoVI/55lVmvr1jdV9Zu
LmqsJt/vY+zkWImpOUUBpGtOcg9e+pKZhiz40CZu5b+TIm24xKfcmw0R9s28uFhVqH9gn2QhHVTA
M3kR3noL2XG5P6p2iuuucSP8w3jcVFjjjK10P0QfOG2zPjky/hIAaAahAiuHddmmuHe8bslSiBj1
r49763B/ZitMz8CSUXRQ/83TUeOQm25aaydaTG0mKph1k83/wOKfveTLAZDsTZHCgk0X6bPbyBVy
EOdhzCZ3nSSA3QIkVC559Y4Db6jVCjqWnBI/gKrgQ6+S4TUGoenc6fJ/+39RNDRnYI9TlY+KPoVd
JSx99/NaRZKzOFINIIuv1j7fV3XeVc8mh+oQeBx8aDknWaRmjY18sGi9e9z8LTp1GqqRAufS8GDT
8QiK23zaMoNZRDYFDd/i7Tup+LyWkFfdErK5X2TfVVzD68EsgUKOJDAgY8rQK2INcSafRHwuKZK1
rPw8vZpHoxaAwVoPU71krafjKVr0HvGhocmKEv1BlVG7dZ81ugQrbaEKEzlVPWnloZW5XbH/ur5Q
QeaI/CGXiY7G8NlbDnXgmG8TFu5qHfC5+fbtRVsk2ZpllZFjX7zRwU3/kdUS5X15m++WujOc9N43
Wk0Klem6uqwvJ1ebp0Hr5PgGWQHK3g0p2zTiGZiFjygR4bu2XJX4TPi5BfeQcY+icp6owjv5ub5d
QVCEDihV24b6rct6RMvceDwnEMer7JW20KkxX1xkY1smBmoVkJx3F12x8MA+U2qeasx4/8RbcUd/
1CzNf+90iAGqIxXsWekaS7AN/AtatjIRhQVZesns61WbnbwJDvAZzkkG1jrYHFx9F2x/BigaoqDz
TljQSf9Kki/p0rRWU3EfA1ZFEcYHjWKV1spwtdAwqmP8xGFL7JAL3ykIBZeCsuX+pDeYGK02SpyA
3liEW2LV63+PL1bLn9v726YH7WYE6Hk+EbdYmDw9Y4+uxW8rxpd2O787TXIEBYt5ltk9K3BQ8CXh
VlPa/eWKSZS13nn/WZ5lymF4oz1+xgd24CYEAxafUdlcemmBo8IG4HeLZ6pjTNczjHhtU4Tx9pJQ
DmV/xbQfsCaDHcymTMEoxqxJPSSMMUzQHqYr7Oh+sd+amSsHVLL1v8Xq2QluZEAYd4+k5CrwsHNR
rPLCOz2oLI9BgGdsbeveJJu/N6vgsmz1HoznzuY1Y+sIWxX6ewuJXVxcKX7m293Ao9AkkeKTpbpw
XB1T/eBQpC69N8htDGiZyn4EBhso5WpZE+Oxrt7Fc+J1fYNcma8WS78r3InTnq87M1+uF7+9bsan
RUHmk/69SSxItcCMOPgkC9ewaNlkRivwEXoMP+VJhFr9k/KqxtI9vOvVYzkNRpsu1CKiMrATR1QG
keg67BhIIaoLc0o5vNuJQHKmINY/OhuFVzpg9YyWEtj/NjE/TF/BMXPujld7spWDFE5G0oBrc6NT
7YJjmTO/kTa8hoymCxGZuBLk9XXIL9fo4qGUYYetaPBZpj6a+LTWzpP0yGSk7hbqY+HMcJbjAa76
Um4tijLkyrH9s7cxBJ9BDiXVHAxHvrjFPPo7Jk8T8EBNAerrci3IsZYTD5uNmkUnPoBOzeQ3x0eE
j6NL/NTEvtIzZoy/2pJNsMDvkVJ/K/Vy76t/jydomRbh+BH0NNmKHKInCUgoGDL0hQbS4hBrlvOl
I88j5k4kfuszFU8JL8JebVf+hfRhydtxri8ZbWp1SNJWsi/az3HQ2niFNMSX9psGquzuB3mQJtIF
InPNlT4VOZGvrQuB0Y6We/cZO+oj5+1dNqGi7Y9G+QoQ2AdG3CRGQkR90vpamsdFx2v/z04SsgA5
3yRmAW4RJBUaVcZLgfHtardQRF8gqLLyy5aGm1lyOOB3p+UnojavBjAZ/+VFzaH+bqUgFgGASdKt
Wp/BiwIPWhuwnjI4jvNWEc2fzepKXScKaSeEYatVZCLaH3Bir7PI/wk088ecOwfi+pM3seNnP7Qq
CH8eakyZmXrXeR+9BeDISRy7LR/lDWxyT13Yq8HWW8nSJ6qahZVxumcvifgFhDz2OJGC1ZTDP1vf
p8OCV3rQuayfo3o3OqaR1kEfZ/3Qmg7J21ElYGLt/S4zvj0zcIk+o74mP0iUDaeX3EG5VavMzPw3
1UXhxuF2+/mdYWY3BhLZQ7V8VztpQJeFznsOB9kAxwu7Br/vXc0p9DboIJqDbePkajIaPar+cp/t
tUg+/oaChgAomd+FpuPu/cskkkdgh2z+CB0ZmdqUysEBJOUI9Yg1QriuTbhT36MBKJ4hWhddKyoh
gnAbBr5bKf0RXAII/CDPvFCp2xrb1ai62J4xncn0i+7zTqgr4Y4sihDjyyWyW345Jild0QCQc+Gc
WEBwRnqVeLePxsPwUdxiCFiRx8zqOYIeN/BAO/wePwz2VFiJuCgJd3cLDaYLQPD9AsEbd07lORMD
dYhf8knaSqUKk/ti5eDnzH4VylbsHMhaC/Kfvcm995mq4bKoTiJRG2o9AAwJYKnkPq/tiF+JAMLY
TZwcr52LXaQLGvXJ0otz1xvB8qfZ5jkjnh5iP/GiHJwzS31EySdmAy3CiIxitYMCi/I/0e7ZcvBB
tijKfnRJHZp5QVrjvPHuDG1MF7OjyTobBm7Ic2GEauCuDLOuZIA8gUN9fC/dnt9xZbkjLE5/9cO4
zeX7LnCdb/EXyRREb+kaRROYZhl4af4v9Ao2xGGL6VoddcDM3UJ4FSHfIwE/6z/e/wF3QqvuBS1W
zGy47DGIktINrrj3gh/QlNqiYrza0igjtXaIgJn7J0aYeqhDSxsuzw6q8MKsWEc4h+4Btnuu+rYQ
gm6JnUwDJ3P3dfmQ/o0/13JL5OxR2T7pF1PU7z2UmWgTCx/LXcTK+hMixQkhmgV5gOFKOrZGElMk
lSE0mze5zXGz/TRcUE4o84d9ZzpKuMJtmDQf2sqyFO8ZOUDH87bNTGckmBQ5+yM1WN0NOkPN0+Oc
OJP1erhlOwgA4cQBIMxax8dHlraUwDlKLtzwORuQLHMQ2MpCC9WcC9C8nbMhRbnCiXLlYeRWH8UX
BjW8otS8M156norGu4H2Uz5b9RCeeiVKB3DuujOjRV2vt/+S5qZ5BSXL61tSHUuruY1hV/91hci1
dszhv5ezbpu9IG8bVnLFu22Nr8dXElG8fnu/05sPXrLq8iHjCaToeIDLuQCNx4ISy6y6KetLkrJ3
LO+vEkx5xVp+VeVWJ2elq99r2qdRHls3DwPT8taQDpMF0AflrqVc/C32liXkwXedjEZiyrITwuQO
Ekr2QQw0NBK9EAejbqUdNzT5+EszNxbZmjYQC95dKUJmvmNrlcrAv7bT4YxzXU/uruLdAC/pKszF
EWmhSNYy8JJdrokkqQW/FFGxS4wpxDxD5cds1xbjo2gtIYtWKjBjS8mQGXz0q541Gu5AEXKy1ozI
Flr+svPvMQg8GFVfM2RY5ay9CSs6t+CVxYLi/RNTXlEkr2jfJECoy2vwu9XOnN3Ce252oIK1suEL
6DbP8TVc2FgrUlHGYAqoMQVe2PfGNofKlR/a8Tx349O8fHJ0Hy6w9LOyOT2ZoQAfLqhVxMIPUbje
nxBXTfH0HXahBeyQpwMpkPGy+jw3pKWqsVYHC+CXnJTcGc3CdcIXCi0Clu2DH5w3pbeMsuBSEMuX
ceKQ0cXtOmXb7AFh5d/Qif/nIAuHla2qpBpru0QsstbvWgb7uVUd3egctevup19drLiMfML0Ha1p
Her0Z3KoeZH77NwMYHs+VWzEpo8qHI2XCMhIYdLc0JNf79ilk1ipb6zb0SzuD/2NOG4jf+wWhkTK
htqmJrEQXsQjypBYQEgxyxYUMOQ4vflByBou5tfzMN3Wwybkk1t4DngeOSfwd4jMUHtIviA7OTJK
tIX+WXcO2BpNm/Aqr5cwi4XlHaivd8Qgo99UtKVqz7QeZQcDt8JFOFFQ8INd/1OwmwQ+Ak9mXU+t
a3EnX1b2+ZTE3TO98EYSflmKlHqVtjWU23bM9OzOHWo71KOGghQXlh9W5Lm+jQyQCFWsRpAQd2bn
y4Tvtl8+oX+p6uYSOocK6a7dkVZZlcKzDZfxnnQCucXShWSJy7yuUnbH0kls0dEdLrdA/jLPnUWT
u+e4PMCJnyKK8AsmIcm4nbTzMhpfpnMZ02wRB8o0qKc6vJZqcq9TzEaSrWUxqt2UsU+xbqqjd+rL
oFejcz3ODCAL8DWXsOvEPrfHKevbbTFqeh6hNO4oSDRC3enJsuwzFHK3xkrbtpG5gr0BEO/nfSrd
viQ/2Jq6pYUadGxwWO0sf6Ec/lyfszi/Q1Kd2SDfwD3M4xHMcO4m2RnnSLP29NYH//1dtzN23fod
yYmfebt+WJGZ1izwFoB0WrVZ1tbKxjbaHIHZU4W3/738wIPIX7tHRkRTKYyVsID2v4PG/2qIFygQ
ZKY/WkO26XsGvQYyPHKJqUndGFE9xDLb2RuqEzK2w4iYguxYYeXtY8AiEqUksLIsVio519ZobvYY
E43oeHn0l1YrcyOgx350MPqAMETdvDVKiQzqog54hkN5F43A/wMJ3QiwVK4rt/WpP/ggFVwjcAIV
NSBsCCsz3hnmFc2cwE4uGeZg3UM/xF1Ct3Hvj2dyBAJzXbeAUFS9XfiPrfvuepD0hBtnOs5ddyl6
/Og1CXEq05/heCVjmPrmLbljKFJMsLo7i5YXdern6hj3CTO/5hkGey29GjfNpgRkS/OBg9hPQCLv
j4neUWbAPBrV9kpSPpKxCdvvMTIXGAqwSV2XIPSP0wcNoYx4sJo1mCHFQEUBXXS3BSyxA17kfdjg
EYR+DlgciClkXAwEp08/A+vFZ2I+B8XD8TbBg0LVwqCp7iqt/9YORNc7DhW/NBbvrOgS6TwfH7Be
aRbXjMNNPfbH3oywNBQz/tlxVywS/em8gdlbRiRIAdkSNT0j2DQD07s6jNnn2nKnY+txLCu1Qlvh
ANFzxY0bM+Tgr9ecFRPAsYfBhGp/OLXIxTpdBDiE4mPgnvRx7P76O3v7CPBO7WxogjyHUEx5gEl1
c6j+GNlvcVxjoi3EZDl2EcI3kf/ulq+EVuYOXouUc1pueXAJ7R7v7lJYvooBl8dUJMqJGUKONC1o
Xu8ZUswiq1GvOUW/9pJXGs+DGJjg8cbgpPoGaxxCys4/WcpBRNLcaG6cEzMc+ajMBL0sLQEBAupO
pl8uShz5gOBAWSFhuQFS/a+qLO/XrQyMoylZTYWNRO5Z/lm5igkTSQtNcsA3G9UAs1/ubedvrnja
Gnin7PLL8RUVRzVJL648eljHEyNWWr7HcF9pMqdKWsonJNKnDT9fUMEWuYSkJlSfpv77H1xmMhCo
eyQAFsK78SrPB4XjOX6UmyxzznmFIzWzscNHuBFYFTVNXSEB3CzZTf8zm4HDsXuwhPHRRj7o8sSQ
ROXYPJPVcxe6IfVWJw1wvDvL6izGEQ3eGx/OpUz3WYRm2891ex5BTwIMVYprAIiAXGd3LzxyIEMh
LfZ/txFrweMdcYWfrEYtaTXc++1SLl9ZrtInwU1QwJji3X4hecLorNvwYCHab4Gz9Qj8nxaZcr1Z
v5nfHGoZ6E2QLaK7k9xQmPKFEIMxujE7G1F7pfKbGWDY0BwLmNbaNpzuerBv1s0PHgTpQvYvxftD
VK8+7DmnV1zkNbcLtd6HUJ1EsgrSLGkftkW6G5A+e/nHCABDK81OwjJUKMTbEidhi6ZTLXZvQ+qm
vBUmGidWU8yvWwBWz6Lndj7NzBPsRpEe1r/4uyTzmYt7syOpkDTsSnPBubm8I5yToI/0lFIJ5mki
0inswN/bTxEiSSo1AK5CQWO/VythDpEUipDmdQ38CwChsuACp2blmdi21q3TnRqDRh5VmXXZ9XNh
PPQ+McNiYMpr3y6g6Yo0Fx6LRKIkJuhRmR/LTRM9B2VIIHOfX0jCHmnJbYzDel6V2vba1nnWbZ2l
pFJB+WtaSbJFBGOtNpNN/zSiUC8pZvnInHI0vRLtOv3KDGllFNrL53KHlGga0a9PoY4lZTNHuPyF
L3lQNmVcUPO9BiuEfJFX8Uj7T7Rd6XRP6LnbWtXZng+SdKXTEYwQIBZiJXE0V/wPPyOm1O7SVr9e
UkodlTaB0Lg0/BqTqR4Vx7SRTzwK5p0T1h7VZGelpE4IwZhbYx/R/MS2+1cc5z8LRzOcQz8fjaLE
CjfehbhMs3AiANChIIjlB8n/S5eJfU4itzNFVZKxUNGYKWf6SEgJHeIQ1nS41e1QCh/qWXM9VMl6
qvdiz+ZMb9GiVxSUSq/a49pHLfc3ELRNS1rU/Y5t+ufs609CY81S52fxeyeEWZNEm6oFY4p9e2ke
pmkLzM1G8mgrgfFbl/8cVyWqCW1UVwX640KzsbJXETjfOUb+iNXR7fjJxOriWth/W0D5f3o3loVm
YLYLUiWzYQ6t4M7Pp1JnAZxFeAWmrAVbqbd1wK3+O40L4/GH2Howojn8Qe4MTf4fzU+99W7Eeg92
zWitNLm8qQJeKN6SD2RtKYlnXlkTYXITFTSkmhTugvdSSQRunDN2i7UsX+KKDbT0X6PoijiUkS3X
9VRAc8bK6WDwHRpSKjJeztoxwSf08nJ5VIJdAYeAVD0kTQZEE0ukUKtgsOSDoThuXinfUa3lre08
NrKv1BldACWlxLkTilx3A96dyrKKFKOF/cyF+3jUIHi+l0CrMkorCBcTBluaLDlM+YAB/kh56NcX
tOCbPokHDz2LDq1hjewfSU6CIFaGw38en/4BpUrK7oZ6awdY4BApFrwYkF4mfwcXwZOidrGZhOyn
inVLM6RS1zfsQxAkba/HiFN71amegg4h46uegLsnxhxluEodJZOMu4yhg5FujY39t3fwFVvLtALg
C5x+DgmmstaKB+dsbeCAiP2yuxlyhutp/qW2xLq524cyS9zrWhzC/H2sKjAMTPMTmXnr63jrkLzU
UrKKR8rFWmBDas9GBC/QuFsPJuo3L3B4cKRfsYYELkc7LkRenELNs81vnJpF0irq1y/lqgi5I1O1
ki+84U8z4/wt17DoWXWpKi4kEa3r20J1X0iY9l3vxBEliEoaF4c68u6Ao8kB0Nstqu2rmVL4eHTk
ZbjXtIJNniqiVAHzlvvieifc1he1QQROQTIMbJDRpvKQt2tsltpHNH9s6/sMIBB5/TNQjNxuEoGm
Vo4QTOn/H8gjthy07QKlCKqf13A4LjtwhY+WBW+aXBRKkg+VVbNE0nqnqKqHuUCUghgnm9acSM0+
ScXGreX46+l8nWdubYmDX0kcHweozrIDj5JmhFKicUm/01aJCHYXyt4y+MBwSYsrFLRCpxrBg3bd
m2nBPe6L19Rr5ACPRlYzRrBANy/ipGuvPGvqUq0hZZtcGz9iFNVcf9KlZ4/tWOeUqTu6am0J2qb3
KGkYQ2EreXv/L822k5p/c4P0QbTYWFYsQV8k+DWlZU45ne2MQsvzBqsptbaIovmw2iXz7F2KUcWw
mX9neMLYa3qqWEr6OaOX59NuhseIoRZ4CdkNW6yVAAgfZlUFUwGKbiwOiAew60bA7xY3jY/5bIx4
2UuykzxK28u4WpZGk4RWsNt7oIhBtQULWrlHHzxd8QP9LC/WiASoppysWMRILOZPnRtmgSFZpuEO
zg4yGHyd+X0Uz9uGcbM6yzAsdtPXmj4sV+q2k5DLSQOE/S9H4SsfR4gjkHCQK+L280brZp9a64J9
r+zZZr/14QoDyTrB8sT/mFy0fqQbsYSDnjShMJPwbJ7EygampbHMcnTUk9KsiboiJKh3Vbex1MQ5
nFJsDucPvuMD0WDtZn8D+Qt9hd4vYS6vyFa+OJ6M6AAMaPt+Tbina46+9+oa4N5+RfH9Ne0RnIYe
FOVgyku+rNtwpR3MyO2m6YmaLYQOPnHurdtfolv2OWYYgHasXVDpzFElpOJ8H9kRvyNLnBOFk5Ax
QD91eS4bG7KCNLngCkYjhCti1uGYIgomOaAtXdpoBFZZg46Dq0JvS8G7RSHDXVe8EHExJO2GYvBS
wmTSPwYd1ELxTfHjE6ks9LVNs8pa4GsWPWlD4+qscJIjcTNCTfAR8Ee6ocbMBJqIKs5+0l0o/szd
XdebCz6uUGWXKdf+wilcrr+t1F5oE4wBxSxGUeXsMfJOXDv5VoymV5M+imMjnKw5rAfRdD1Oi74h
TKJxwuRbsKmn6ju8VWfGH1Cmx69uNdC2IWUy3lRXU+mpx6Y6WdOT+LQSGhl5HM/pPQ22G3KK0H1b
v/S0SLyZtguDOD5/HXlufMlU4nl0mh0QljFsrnH36/UuqmYHjKnA4MRHzaC9ZT65w7G5xUa6yGYc
HFywVffCDIJIiTQmohZ7IowRK46K4vlSB1xioKs/4wMmMytx4mB+fqaTN476lyZ7eN8Ck7fq6COm
jgX7WTCSMaJ7hcTQ6V7lLUs4/clBYrfr9H27d5IHL6aDcRVM/GM/OpxuNOebAjIiMx8+KvUJusKS
rGUtXBnOwNH795LqtwRhFZ9XwcESI7SJmPH1jYtrmopXG6/8rBjQ56+7B3FLoBHG9RJvrOad8SUX
I+X/NM7SoflQete+zOSB/AmmgYkxtUPN5AC3P2MxdqWKvOyGIyG4fgzV4zC5/K90STMdOuePjYfd
CbxTOwapDYl+v2cqbtbrqDqiYoCVPCiQlfFwhhe6s3lArPNa68gfebLSsmhtNr4DdVOdkdT1Qfp1
4BlIgWMufDTtZQTxOGgWZWyEpEZ4vP/a9ZS3i1kxSmWjaBUMONSsmTB4UHKgP7sd+uDf5wNflJwA
rGB2b7FQQw1NOVpyE6ABq92yvheh2H9UkbPYPtK3/WJDFplEEaQHVvNX8G+bwxsmgGXhfRU4uvir
8pAPrbfmoXKV4spnaLs+G77Du+VDrZFssa/917teB3MWJxdAaxHKJTi6tas0vCitP05mUAXpwI7K
WBJTo/1YcFEGe6YUrkbMnUfDcOEXbp7vvTqmddWFEG5hjNb3ltJ0AfEaTAFUrH9O89S/mchNpMCF
slYq9x8TtP+J5VszAVHZAQgUM6hFCZmXMNTGujTC6Lhth7c0myoq3HYibR5iHxc6VvKD/BfhtnKP
kYrNqWsrKqejH9E0/uyyiNBEHIjpH8XaCj42Haeko+gQziBumGUrdG84ox/x7p//LE6UOS5ciGRy
RuEozujRQvXjKLYA3KQOvlA0zHBfqfvzduQb37kx9jtjqxDOdqikxNE7oKcSDnVHyYVCXij11weH
w0T1YLik9nA2pylrq0Fwqftzju/RB29fV8usFUBwoGgGNmKvLQxmktlC95rDBgGse0iKiuPvibXf
gUw1qz+6gTsh9Ke9qlMNS9iEx5i/5uFxz63frertuHJJ+/c0JN8Z2NXSisYNot4QKUwfzLZguaIL
UQXF/BXDo307znqcCQi8Yr1pBIhKwSMpZNktRFTNZ2FMCwGoW0h0vAIAiHGTZFZFgGgrwUOGf4oK
VONYxbr3yU5I2+TpHJeqMZWKWz4ODFPTJNuqEcukSG694pDe9pxvxySysT9EiRiHISG1CkqEaOSB
/7SgKyohuYkSjgbfW9Mce908KLGQ4SkUBJhxCF8fAb/0Aw9VsfvEkGPuTH9R++QuzaTvDcq5xD7N
IfJatju4kqNpgVPGqZGqQPNlF8Z2GZ0BnefcY8C6AmiXiu0FEyV866cEc8psbV16yZzpwHRr7eHH
tHAfjK94+6bilqqaeZT0Xx1Stf2aBbLT4mRDSMxepc2vxCAelC7k9UD3wj/Yj8f4ujZ4/Osze69c
MrY2vQVETGYUXJAstIIKgSa+RI68Ncy203o8zgpb2TRKj6yZr1TJ4/nwXIaKj3VIaOm/wA6klsmx
s6S6cdaoEmVz8MgPfsEbJNQYvGE53uDn7FbaMAkH6RwPKgp0/y7UrD93gngcUN0dEzFsJ/1/w7Be
4lhpv0mQqUzTnU5nM/oizFunY9rdOMsd3UkHTsQwKgjthhMTUi1mE9k4mc24RSuoHfzcj+PpswEX
fQfL2D98feHUOaf9FWqDkFomiA8xXJwp/QDUmk3LnZjHS4A9tjHMj+UQEfYAaNltwttvBnaW5yWr
7oEt6xEBTo/VSIhpeAHvH/IsZ8hT0IMwB/T5wlL4fmqUTn1bmGRrnoNAt60iUV+TaKHHJbIuBvJd
P9G+SiBaADiOwq0s3zCC01UGhwPnNRxSnyATBVGPbf7Kyf4Ofp/UMP1DiXwsjDVbYUXytPNr6nZ9
GcOnG9njb67GXr8tjAer5ILf8lh9pHScV3c3NSUPQA0x7T2AQUsbpNT9agLVeiYN5GMPN4oNF7CA
VzL8+z0jEDd1+smXKOHAV3E7EDxD1JeAheNsCw8OX+G2qAOPqePJFhC7lQz3zdPd8G8Ce0QM6oVA
q6UQJrD7uvJ/q3UYIqY+FG8HgCoChqacQI3OV4soAdpnWQDe+AVPZ4TcKbZ2LHxrCbzZ4xgXLhsA
ZvtBslwHd925fBhxOpT3Y/ThNVvIxTgx5mNrhoj5Dzn+EmeVZk7He3YnU6mvMRmT+8kzN1MF0d37
c3cmv9gjtW8P3EMjGs+IhVnC/XkgY9eyQjp/YHDfvQaU0o2p1h7SRhKSTUgNFAWEzlrssvdcCWw/
rMkWU2l+iJ/aQGt98VZx7V6+2RcBxsq7MCfL5edz3etOP7QTjjk4DpHEdqbNjiJGgsW4NHxmn3Q2
xaeWKXjdLoaC+9gHygyMcGDMv7mRZYKvYvML2b/cyfeP2YROz8NxJWG/ucL2sk8lI+LBY/Iv6+Pw
hYyUgwdS1DZ7OUwsVanvCJ5BfSA15pi09wKBcoEJWd1wN787bptyQJNd3nnQiFQfOHuxJJ87mOF0
U83EYuIgAMFzu/qvUGsi5ezKWAkJZ/8FaKG2TiUOj9Y1HnuslpBUCecMrfJHLgysW8zMvg88kDEx
sY5lW2acwS1zfZF7eOjxwer6VtSTg0aOXOAtEFPvu7jXIwKPrEofKVQdto2Ux3daTy9p/iYhshwZ
hj+i2ibf9Zm5khq/d/dL32+Tu/efMjzRcV+XI8PkjcHNUuwaD8SVY2OvAupiw1eO5z6K8/GuKiZ+
9N9/tqQAiEdcInEAGyq6mhAhYWjmmvKHKaOT8udZmXq1BdusvwZwyejKGfmK6lKsv07IvdLK8CJE
wlvKzyHoBa3gSgeu+RIcUGw6Hskfz/S0SXzyPcUcylGxqm9wvV0PSqqWmVzrknZr0vOxzi+T4Pdh
x8T3IXOZqF8A6yGlFkVfflbpa8VWxzvivzA3gqp1YKjkoGR6vIwlFGzSU1Kix0tNY98mRU0n7XkX
8kzi91mcFoErZ47Fe6kV7DlRsnPTwhGlO7sp2RIIiCDXD6g3GTY/RodduNmlUM9GcCAjzHuGKTNx
/0VSSyxZjqk1MBYGujEM1ZtOQ+VTyNK3Rri1hX+p36r4f1TnoekLjGKr1NuMEUWfNv7p0uvbtIdh
Ie7AWLZ6eatnQWV8bEeoE3JlVC7iWyrszVlEbAUDNpxC5T0o6guSoyxQCnUtOQcfzXlSCDKgj0w4
hzjDe8h6aiudl4gK1w+y6BJRJMdHfK4riZP5FKnvJrsCMDDgL+B13inlC7uMrpFBJvqPiKwUVI/B
C7mdcTnE81zowgMiVUMUmd16qe3uytm5EkGDYVe+O5anrKsK07H1Ea4CPApZjkOYjmDELXggqghk
ZMv1a99MMyz+t+HjSWgnXXP5fBnNULW2zD6vrqkogeTxQazZomAlq1co9PRZSmCjtCePSWKDSafX
CvKxJbmIrHor7JOPE7MeVB+yAfli9vOFKgYaMp46e0ayvBD+u7gtNSW7xaim9G3qnmJLGP5lCxBV
CWtb6CyZ7W0G3ktg8L8f7XJqjdZ8wms/KscjRivS+DImiL2pW12Z1/65yge7KpWfffnotMmqhqW/
mazxQXlJL8wOOnigRENcKe5sYF6PI/UuFBBUM7iIkdctKSvVDjNo/JrpxDgZluEiP0zo8p9NI45m
ramtqlKOP1lSPmSk+o8PafBn2Kzphkiz8O7w6ji8S8+t/D4vKOjRKZHrGu4b5cG60B7B2SfrPmhx
GiPCm/UN8Hh69ef6ni22yoeIBbKmJgSyA93NTGYRHcEtIEf9Ka7mK3SlVzmjd8dQW4aE1d7Y3nUn
LJg0ybMHH52eyvAaLGhS0OOhy5Xi1mnU+T5dfuYVyb1SRQ6KmPVlo5pq6MX7s6fmVZ+anKWUTwnA
tiwg4bJsvQll1ko41vxYAlpHiTvVmnyW6AHew70p0cvdmlZhln+OywxqpNvqhdrP78JK22jE6qR9
jVue2fiSy9fWXSsS7Qah+UYGTS2enx9VzrCdtXKKLdX2vRTjcULE78Y53Ks1HE+J1xhlaDjYpVG3
t+PjZ5hNtT09DaaPp6mJA317D2rFnrJRM8OWW+VZRkU3tDRgmeAah3kez1CBC+fOUpbpP5DWaWcp
mFeWtvaH9445aCcb+zQFNSGZ3XovwJpfgl2htcS2uN3UVjzgy5z8zNHoiIFDHqnlFpOcynVdrw3N
vpqJYJAkPDa9UJnWpTEon6sSf/ZY5Ppl70HOC8ZLt9x6tAUsi3fGov7GOEgK3EfZkaySWLHzXPwt
cG9ATIFKy+K+tmRKsIYu0exK0NVNxV51R8cn33X04hr1RT4qh8+RQIbl/bTFg3PpDFia2A+lat1n
N7GHvNB5BU/5B8ts4LMpb7SXU3XhNsOEuQeNmrTkn0K0a8xEn9z7T4gTh9RxrhybLf30vf//aRm/
Mb0NuTqbK+hndsvqlvGUUEgk8CAXin6KeMtcefbaA0mP68z9vNdFvOsRXaq5by0lr06PksgfbAgP
L7ClFodXj9LSP2m3mVIOzhtKDP0TTZAd8sEzhvxEuiVQD/FHKsP7/TXkFKwj6KHXDOVzosR1OO2p
VizkwuZ01r0NRSA1kkEkBti1vWFm3s6xmlUup63x9ADHENtHrlJ+mV4PO2etNZ465W8zVgB0YiRM
b7XwjWxiwdGlPBtZoDfArQJeYn+GmBVbsTX3Dt3wj52aHnw52u4xfc+oRb0l+GTdjI/cgzYKmkl9
uuAgzq5dQgcz4lCbFrUhc9RR4bcwnR5h0ASwg8VrkvqH3NnuILn8N9us5dBP8/GXcsPblYVWxTd0
CQ4p7iH7nc0rxJcR1XXIHEh5vpiFoftUR1gpgGoLMbWzWF4ELWo50oFclSOjZEVC/g+h3v3vOdl7
Jts/X2x2t0WK8Asax4JC0pdr+9Ix2OWMTXXk9+oU+5mfYqTc/9Z++Y95aoJL0I3rZ9yT2xuI+kdj
jEXFZpObRczWzdpAznigLxor1J0EiZ+7ljTYF3dQV9AlCl27/pvL0jjmKSxZse4s/zMrfAkAs4uE
EHRQhjLGidNtqZwBa2P54gleTrQPk/hz10EIWp/R8WUyeqXazm0CxAUe/1t9AfnbaubES+F2BR1u
kPtNRCgYjdoafn9saM2Gujgn1QhlWHcHXry/tLE9s7PR/NuD32aBC9/5WbV1Fmm55lsUPaHDrlV2
qrUPZxa5kVg9OF6VCEIvCtJiRsYJeMXAtOIL49xRfCG+Q3Ir9ymuDgT1l4EgT/DUynFqAS+GwhPe
ounj5aZ9Zf8dMkPyAHwMx2BKNfsBZOGIlydS4oRGlsTsQ5L0kDM8gR/HXKnMaZT+IJDslI+kWNVJ
PL72F9s+yb81ALGgAOT506b6t9Hn/iHPcucMZWC6IfN5YkGFVKWmFr6WUkWOEtij5mttUS/IdYy+
hC55TaspmJDJ8A5/fbgmnC6ouqJ6R/KkG7HkmJDGMRx3fE6lf3PM0ulE3qYxddmlD5oXQJFRDDDF
j8i3+EpWU2fW4bXwIdbJp7GiKxiDEdQ6MWMsSWmvP+tCxDjW+zNQaSGUezL5j09OvETc692HDgbz
59UOt27xcR1EEbF4SMH/VmdfxIFNntO952SEUzwkr3Q0r1+oemoFt3FlY/g4PdiZUMb6/hnfLO3g
UdEWm4Vw2abmZ2ua0PWMRRBbHv+iifa4ErerzlvfmpRULAaxlBc3DP2oMi/B6rGtXhXQ9npG8dMF
9BAtyDloR1EoU6XhMIKpFdj9E3cfEQeO1W4Rq4xnuBm59e1p7y2sHD0Ij3J5l408rUoXLIWM8528
7jUgMazdDHlH/nfkU0Zvw8PTYlwNOQ8rPOseE1ewvoZ09ORVvUmTQC/om6YhKeoI2ITbbegTEiZR
2P8uE5n35fAYr22Ttpwe9tJ62nSjvj8WKjqoVQGuROyDVTHKSqCS9nWFNqQuF4rNlZHR0aNL57EV
4viQd72hpDx3xrBIXgV9V3TLbhxY1R2QV+4DPr/UA1IG2EfuUpBd68K0ofXTwsVEvR9X/Kmfvwry
/2ypn4cFpxGtEwqsvCFPRuh37MqefxOtzChyIFRpudP9yJxBmmmrqO8C5ywvWQfN64R0uGEbIc/0
S4LRjIpJpHmfEmOcEOKHgrWMwkiK9phsAZiZUGYEc4La2s8S1dCgiaGCVWLt/RrNKsSydskE8lxM
f1DGlLw37H8nAHaEPG+g2x/vkoHylC+lhUGRJgtay7Ynx3PKvysY/dlcp2dJSZ2LnC0Ea4jSRrqS
sEsOu6UtD+wO9EZwahBEHyr9girLMaOgJNZShNS6FZlGacV3A3kvQE8nomvTE2sOZOkrC3dmich3
iZxgU2gonMFMS6NRnU/fpxsUXFmsKbrx3aqhuzMaywscDPXtcrmsAik7meRYKgYc6B9uqW6+fB1c
rQd0mEDxLwlsk5NsQJqyh+cJa90hC2Kz7t0GUhrGApFAFtgM0dFkYK3jvBw8/uiyD37TIiFyVs3E
oB/mAGdCEvjrmQYlvzmzb3c7MzNP0lyX+LYNyhHc8iDbAZuXDfZgjN+qJf4ammY7oloCtKuIswl5
+BF6dIvuV5F5D3Y5FgzhoLmgUMQ+H+AY5OYaSmeHM19m77XWSKFSxTDhT2rgwJEU7M/3oiwU9Ym0
ydWCbErlxXGF+Hf4/leE5A1p1GE95XOFH9O0FYhueCW8NF8WyeHxO8xUpCxN1jGyDA4F85PlVgrP
geO9nqnDD/d8A5o0vJs176418okyP1tj6sfjd+hbqM09JM1FjlaYoRMYGmb4B3zhu+82hvJOXaju
YvKucjuApo/OL1724Vce6yJc2NnswFPzFJq+D/Vd9zJcl3Xf4N4kCciEK/KrSLS09ejFxOiX8OrB
Dr715qeGtFqg+UnUtZ9ye3IPw1c+quu1MeWe46Fbk/MWv/1xAmnBRqMZ/Ll1OsteBgfM3dsI3z8s
NottaoFbALNxUOBNPyhSBFLnqdhSpiDUxcncKgYvck4UJVQSy57QMr1aBcprg0UEYKWWgOg0Ijy3
/cPR52KOVRJp2q1SPAFT04sSxaZLRUO0ENJTK4ai83/7GBcdyJSYeHszb2LdTodDm2dEwjifFZ5N
h3mUtHGO1Q7EUoyBELXv78uvQRRqov9MGOQHwXAbBZOQXQMPwXWkco5g+amHJm4sXIHts/Tvb4nQ
UzZLyCm/jVz4SQgtTfR7FWGZT5Eo4AL99q5mbBMNtXQpq+zo5H9kRnzAgyuShDkSDwOLAodZUOEL
BTEafxCjMjhjJIyEIGIRHLY/4QgmpNIYFN3QwEg+pMpoaVFCMMS/YoTp/hy1QIu8LMZyDXCSxoko
LX8+tSO4THk526Dgzqoi8F45Lgy+3Zd9zlafPedCpoedUEUlvupaVohTPIdJ6ANUQewQwHYyfjje
kwgPkzF2l2ogqcnIQAMOcGlg91uBsrfMQUzF2hY7N/crns2XHfAMN2jbmPHi4hwg8QszIbwK+f8c
OMTqOh8GCGOHUaVZn8bksGwRhOJFq/4O+clG3LQKql3CMHsYWWkNX3zugtw3TPzD6ELH6hfApHfG
JlXjebilPZk/m9S9WYvYJFwpGxZNTHsKcwGgIbF3P/qyXxvVksq5lnjjrPhWtTbToXGI3IwKYBxs
8O/iUvjzEPrn5bsrd7h7wQTLb2xnK8O+Yr/zFPrb33iq+VEFWgeSSzo78ESKlpEqbDfFUiFn6ve9
z2LE9XDjTcB5LX3vM5KcznJo/enKJjeGjQgT6T7FcjfFyqClp0SutWd8Mcnu04EyWoHRGlpWVeaq
FcM2nsRuFH78MALfgMHR9Dkuw7P2raYcUzKP9LV4q+hJmx/w85Jc3ZW8vMzdyrgp4P12I2G9u9kZ
ELdz+5Yohjimbf41Pe6kuYlwHOgt5qbRlMXs2sj/Y3zhOECDK9EQr5yF619UxzMqYAl5dCtK1aWY
vfZnMvRzqlCsMhMx550LpwYX8HLErxRt7YIHduS5HuQYOHeCV0yKj7Kit3pY8Fohg9CJ+VNLfZ9+
8a6lCg+KE9Bf44GF45XZbsePxhi0xV/2ntNXRLicloJ64s717trMTLKvDcHKK/8SA/iJw1ic/2WX
MygJFl4PPBD3fqbm9iCeDQYU+GPllvbjKduG/kfReM0X/GamR6g4+XIVpaTiqm6f3tJiT0YoHNVJ
/MWr3InGWmQsX5E3AX5t/aQ9EvvyZ0Rv85cEdqy0uxM9TJFjkjrm9A5AoOcwd3tPnHspTaMmzR4S
l81wvG8w51Lr94xjw/e1SPZDYk3JOYiezhw++F1LM4yvNu2t29dtP/kG3YohWSaWT8hVVlxsZBHl
yxJHwq4ghSxBvBRTl4u4hEoq2zXSNq/zaAceTXTr5FCiIluNeHwlwfs2UvNxnEd4N6lidDo34XoC
PAEVwoO+6n/OGAuT/a5OxpNqx0rZdlzzyWdlhjJR/70QCZIJVHjYAJVqjXd1gNa8G7DF0nWwdCOy
UB2AYUZp7XEo3XOeCt/4VGn923ww+BjN6kPSWTwtD9yTwgqFP6W+0NN90xC2rmhKYr/4QXMGDjx0
VF1FIYEC7Ju+vnXnaV8vUTRcFxnJffMljcPFomMebFWlqcOinrvtoRzRmfscuCSHuJj8vJ7R8puG
h6XWePpvgngYpGhXz7dnBrxRAgoX5h+FjM+fPCZv02cH6OQ36ioz+tx61rqu5pN5gyMwUqVxozEP
foamtuO+3CkUIHz/UjY2Lln8WpTG3UN4A1zsYbHIRp7oMocAOnZnxY9ssAkk6XGpf25RGm4g2Ldi
N08kggp2FV5waDWuja0mB3te50Y7LrWgHz8cQbaZSSw9FgLMLgpBLXmdSdj0fr4U7G36gsgHnjn0
MhJYlwZYMZWDUbrsu/ZsQZshEAiOSo0qh7PPHjql3bGiGX7RqNFFUng2fdUsO06pEkW3zpOlhn7W
ZXragc4ayJpTM/p8LfbVJE/4ma7G6DXAM5zyfxiUhlYtwgMSH8Q97EoLha536WEAM7NXzkZH+I8d
2/WemLNTell4QE2IAo5ghRVArmZcAGjEF6CO8oHQ9tobBfVS8z/orlGpe1CLeGkYzU7RM8gRSlWb
ZJvdWycNtgd9QjKgGiPywcbHzN3exBs2aqCSTNVVBbBHy+n1fMcyygrW+NWvWzSQj96Y90f7YRU1
WvzhrNNB91zuYvV9tUQm3cy7GaZn3iI0FVp5LAYaPuvK0irlgHia1JtXEptcJqGBkYiJf78rgCj1
AhdM/9qOPZ87Qza421D0WZn13DzAZhvtUNETV3+WtCSD2/ZyCfmY8pL/d+R5I1q4RRvwfijlliVD
wleNznxWC+eW7ybAwW7zl3vYihrRwpCs6mn5DJCh3FH2H1Bv1ExrG+xmv5lvkYQm/FoNmLdW5VUn
EGS0XIy5EE3GiORxXMDTRjjqkq7+HPEgMLAoZhiOumxebwVkgfFRI0t+h7aEKIg8YhErmVrwZfVg
I57/gSKRQ4tAjQPK94jJVSD9wYduTldxWnwZVWE5IpNNyf4eD1k/D3QBvIu/IbO8712WZK0r8xBt
/OTb2oe6Ou87v3FFberT1zOp4od8PvEjGpYCyASh5ePMKc8Yo0pZKhTUC0vDxnfcd7kXr9o6u5TI
vGepVPClS317Q3MG60JkkjAg0rNrKgDQWH5Tr8qIo3kfy7VYxDiopurIEZnQtiiQNfNxRWn33YJS
9DbwlfQPv+q9aJ3J2JY2xkJeihmLCd3r3vrM53GnTNYKDRdFL7YLsfqYz082tyjBPK0xZgTgvLcF
msr0T0EPviMO2S7LOJUZfiSePl4pfloVYcUvBGzXP+QLVKu4OWNHCdZysM8JmK4eCKQRQiLMmtEL
u6rnke2LFN/lC1gqynKhxeHF0eP5M4noZR1ib2jZkAjJlDGoONdEMSkK9nVpevx7M3Pv0EW4sadX
B4kes+5Kc63nxE64aevc+GiJd2EbpID2bBwTiaz6NdPNSxUy6R2Vh0Oj/VB9vo2v+ZYwO1lKQk4l
TpLJgJ/GL0tuQ33bgjSOHf2uLaqtzgfPyYkZtaSVPIEscIqXo0DsmQsSZO0M9Np9oPkD3E50EQuc
N9S9DQS3UQiBw0xg0rZL6sSHJ+3ZqRgTjUuzfyHibcbz8Ibv4A91VS6IPx+LHjFeTlSztau3f0BE
r7Fok7dycyNQoNS9hn3dn+/+IB4AYSszdtddeaut/0+jL8Q8Nsjba2wj/XavblrvznR5a72xGasx
J5tp4NV99ZUq9Hf135TtTpOZIMrsb7ktcumNr1SrdPxeMyRRnp59uOTVc3uVQmkbKKGTaus4VInD
ocEBYcDLS6tbfzwN19fbhY97tIUWz5/J9QF+RAq+nmbpCV9K+HYxqCiFh3wzCofMg0El2bk5ny2W
rSgR7LQYiZwe4bMkGtOWmsgYEaxlU3wWH9Wrg1q2rDUXpKS+pz8jJoMzhRDA6DNPbL4dE1qQBq2l
/mtKHxJaa5St5J8vBh7ImOwseVq5UsEUf3zTixJouQ3i99ZB7aRppQZCntzyaqA7a3RN2BqQYNKL
jIFIct1NuC6RXMcMMQTxNm0ODIxzu16Ezw9H47PExXbDq/VX1VEqk8zk9un08+utzps9DzqUkrxI
XKuJCVUcCYznIPYL70E/fRn6HbHKJFaz+x5FpKJu5KuPHf6gqboMvovmUeO+Gf560TMCGFzuoCzM
FPvrh7uyyviFNVZjFiVqko3AjNqxfKIJna2O77ei+p9GinQwKiNde7TBiKrHfVKWp8u/VA0lu/+3
kWn4xleYTFhxlTz1ADhaD93hVPB7GMrwyhOTdXBUG9ZfbRGc4XjLoaQLyuvvXHUWp7xWmnXh1EeE
ItGqV9UbJOJesQcxHiC7iKzRuk9KEz9vwQwSj5qlS0kNTKRbJlrinBurR4Y2o4CEJ/kM8kvcqiPK
incmwUxMzvo+6rv13Oy2y9BbMQfaHtOxhTk8gpbZNnbFf6iLgla3JHJMUABFvffmHY0WfWHPj477
8FyVnkmaLqGsQ5G+9WQ1s/4eIh0Okz9sUm0z3Tg0W/i5c2jiSrslKIbL9kdlYhBFWRODICEFHbfs
UlSmpMEawpQ8MfR2WKvbQOPC+7oTsrE0jhS4HnxpFfBYriR2Le6FrRQm6IBKwBUjtMW36IwexQsK
VMCAxr2JBorKCLDKLw8udo2JHiHTW/q6j0MEKR7unQ7V+Z4ma4nM+xuiEznnCqfsv80GjGZ73D4m
YLJ8EWLktHRgXUCebFGRuUAXOs5/FO71toVZ5XEk5/IxTyuOB5gRNvYCILwvUJj3fq4Pz/dkw3UF
Znos0rs8EYa7p7isbXbEILmMMvlMOQ71Zb8meO5KFheHHITC3ksDq0cWIX8bqyWTmE09+hwT96GP
+01saK/5Lqu9o11q9XaGxRmaGtalEKSo27neonjPaXUS+3pe6hv57yY/TlQc00Q/wtdWu/6WHPKo
j0CdbLNCybl3euvhw5GX4uOLI3GbfIwKAhobBX5pp1STzUIW2yuuOTipp3n1R8SNrxhyoOht3o3K
lVRleKv8zbuoA2ALa9CAMRWwbQRye5haggg6458rC6veWdo/yEza/QD8YRJb658F8wVExInK7L15
7i4e8GTQTtsqY+p0GP+M80S5AQwEvFH/QRcAQVZb6iUQU/uMER09TinljBGMNHQ2osqgaRCwQZ1G
PMbc1XvYQ9SUnzcvpC9cMRmLAOc8OSaxQa7PIz+PPcGfYM4Vt+2sLs5gi/fgu/PNLzhGEJb9tXFT
UG4GtWeLPCum10RZyxqLGuhNpb+SACBsN2+VS+lSbNaMaNogdkuX9//EBtHbjAteDvF+gLDSvQNq
3oU6WDWTuKvZjylad4ZxRHnnIrV3bN0oPJAYP8rbW0NMYFPlro5AtrgctVKgm+8czxJaPsyI5Qrk
td/zwDG3sVvAZxuLQZYBleYAEwsppGmJYO9I2K+GO6bFyX9zLO2K25aelXBsi+IUtYDs5SK6RbVd
ug6GzGPC8Vi6DqBuKRrEgsDZfJRxrHqj06xaE6l3t/lirG71qJqSdvPBx7CqJtA9MqN6mPkq1jpZ
gy60mty2XNzK5vWSOCHzxhV7BK7OQI2tPutmF7W4741glz0PFF6fR7xseT8vEOiw/eIQd95c1Kw5
+0gN08DcqRWH0248XsO4xdhr2vdtmQCaAugT/mTNtQ1g/uQNCrbA2lPR453NQvyHLnx2rLIimRZ3
YGMYjw6gP9VhWg7BpdL5YMlwglMRI+u7Sxh+E6B06vMzR/RgLhfM2upSDX9uynas0wvxUxsD56zH
hPl0spJ3Ljb/Iac3BPNOKQhWIqXW7Xzum2BSFOoPHZfnNHEphMcpr6zwERktavbDBDw5++79K+1e
AWS8unK6ndrcIIrmYGxlCzegwib4yaobHiEpv7gygLpx6lZq9cZjak9tkOdwkadCo4viEt0XE/8V
fy9BVramUu4Mn74hklXfb5mgM7Yy0DRAmem2dKQB2agsFBciFO21UdGWBglVEKpa+0LIdVVcp0Aj
+V67YY3V4JrgZbf13/EMMXbO/6h1L7ElhAPY58AG8ldMF3PuEXUydIk5Iw0SgZhiMXHWsmaIp9pf
iRfETsece4jX7C2GY+16b8wpnRJcRxdVv8NcucckYcwV/k3poo/FJ/evpkzqLMQ5FnrxHaM2INJR
cjynkWvy4DnUy0ELwih/5Peta1roAKUtvB1X19rLyRiMlg1VZkt/xiAIn5OyexzDIVCWKRxYr6sz
cTkE8e8ScxZ0YVxzBgMDe+tgKDytm/NDjTz1Zwj+mv/nXOPdUk/z+8cxSH7MU2V+tH+rqnf/KIZX
xGuRyXGYItkTv8fROiKMggv2HgaHHpbAnFONwp0tGq573wFG41C6QWkg32vD34bzg81LFCD1FjXS
pEHoJT4II9qOYoVAJyArAth2JC55/9UVoNQ64se6ftuP05P9S/0IGhze23bDADOFQMhEwxUe7Ptm
07e+4/4kYEY9vxe5wnC6pzJt+WcQaSqLkJAyNvnXsJPJWqZbYA8c2YomI1ZLggTydejX50oTlkSU
QSUUwl2dp6Ak13ppy/83nS5x0/VR2mVVeotCx4qdYUIxhwFvUZufFugtnGng2ozsQPHLrfQRXF4g
VsLn3G51xfcOLYNamHCSYzVSIgpqlbz5ppLGgHKJxVdb0Pa15y3GicrZYGkpkKruDMtgLLEq33Jb
MU+Vp/wRo9nuYbXSjm0o087L7pt2kS8ZAI0JvVi3nuLgWj7GHghDR8CrDIYJdoENGrkUnKbWiKAd
42M+Lj+4rHIGk07101Nx8h16l3pXmfXuuCSMn5ADdw02yv2ye+bmzTEk775vFXzdPFPnfvSsDOjA
KqeVhI7avLQpYSAHgH0a+Mhvr9XrYCzo7Y1kINjHiOqunbM9ggw5ejDHMSgmAq9IbDuW6LHV9tU1
S0Dzjz58Z3bWxYfMJV0DQjMKIhhfQN5n4tqz+etLus9xrfuwNioM5GQEfTGSXPigL64TS0i4+Vha
D3AGCdpKM9VAfqCBjiqu859s9j7+vleOEPDg5CHU/jwgbp/fpH/fnTzxKslk0m8D+4cTK7HpnxXB
RDED/4Une5Gy2dH0capxas0dZqNXuEj01G4MJ8gBsVxOE97eXimcsWxluVVDCRU+hT85tkpCU4qC
zoSDROWJ7EONVaoJGfLZmy97k0DugY7QKdbv8pKbYUgU3CWPuf8DN6u87vQw9Ly0RnkS+kzm3nRk
/gRQNthw1JTfAZA0QzzlCCAzHIWg8FlhiFtQJ+9RPi/cTifyDkYko8XJ/3jDUEdV9jjskY/eiMcU
ArkR5/sdsXP2SgZiZjkD+HPOsPycud5rVwYOy4QrFmEA6W5SPd2XnS2h2XNHxrL9KVmli7uIGvb7
dJvuHmoOzq1mJIN0rcFaQSBstbQa4G+bsuATkPRI36PvycCdKmcgjGJCkAFr31gdPJhQGkzuCQa4
3Af1t2hqaK3+I3laCojNqR+oeklCyBygwwr1Zl7MJSonJ7dlbJkt/ZiEbJ9P2DgDOUv9E0YrPqTJ
Fmk36/5MMbvOVg3Zso/BUkM8nbmkEepgzks98IlVWRQAQhF+7BaHQM8/rWdZT53NfG0DZtrp28eh
blLLQJNBgZw0NiR8iNHVD99QjkTNoXAn2xjPcxGStr1MrDWz4cPn7W1tSUdDEmPgL/5HccgiZD/D
ZKCs7UCdbljonGRe3MHYVwmR5O5IwUoX/PKsTgDodIucGY/u3R4sBC10sD6E8avqfSGaE+O4QN9A
o4DKTE/ziB+lUwBAEpsxdIelIan2vQ6gbm+0NaSgSj83ptYShPis5qviic5wquiKINp7Kk6wREIp
mjKX7EfjeKuXaklj8lUfO+fF0RCmb/IOJmi3ksYPA/GHFQR+ls1nKE3wDXkizML9uUqwoRIG4cuY
eF+6T01zTqIIcNN1ylASI3Ap2wrGn2qlUEE4ejrCpWaaD3IyZGal9Mik5RQEsjaMFkQOyzUzXthz
JP8LKkcQtMi7ueHwWiPupS97CRk9r6MgTj8ujhX0emcJNxM9B0Guc1ixRTqZ6vCf2nLUuYxmO2Vz
63M6wX62zuj8Dqg6IfC2balEYQHFDKuIOC779VG7lZsFjsk9FrvUJJQAAQ6l6YQKaQrh0V04O9Ex
b3vIdqP1WcO8ueez+DyQKS9InjA5HK+U/LO86THwmOzid0vfm2MDqXUVvQLvdwMI9TVGHJGl8jSI
DNGM+zbGogxcV81ntDDWP5XiLEs4jNlet/gj8l8RRu9sQRAapCht7wV3sBP0aM573F3zqOKkST9D
PeKX5kTA3+haf/0+uX+53jhoGPYkf5+73WVEIf2DzywhepLHNfrWd7VxF1R05GTo2STRQO++j5E9
dPb6plHDbtzSlujUsMHjryFs2qgJrGWTK+j2GH4Sz7hUobu8SX1QP8BpUzE22XpjbeOy3fa+8aA4
ec2AMWcEjFXh04gXTv0gA9o+H7AGcsxUPcpTyjQl/zm1+ZUowSLgJp1jsO3dejn+YiVox1+FHVYW
dvz8XM7JNqHKEp2T5+87EqtTpHI2fk7UvShk4ymBuRshCrb2zVCfNIYYehToIa4tjOe0ZBuhfPpc
5MYMP0s8hJANybBirNVJbPI+6cgudFVucGnUML95sGmSRxamXlvdc0kB2PHdz9r8ceyo952Huted
xXlPfb4M756qBGMcueXUKPs9xIodIz6kpfFclv9sC7WymbOZxznp9jRwfmT5TevgWsQj8P8KIlWf
222DF6uPGKjRZbONe8WE9ojk6yYhR7D3jkN38CIBwjstVjRj9/J99QqZVw0GpiPJdTG4TzuSqVRl
1p8XcCHQm1FRYubblFPV/4tG9+msLf931fuL9vtKuxjop+GzJdELXXf4mwGxClM+5siLom8g9U2w
uOZAxQ4xmfwSJvZdZjqL1+QrsvtrSe2wWFMQcJxfOjuIGo1Y10/fG1ncHIAwgtCWF+kra9KhOSAC
stHPCyIR7Wqa3laA6Xi4RDltnOtp8uffI4GtN7OI6cGJ91ho/xV+vV8zhvmvCPXdL+Vz3kySoLRu
aIKogoap6ZBOVVz2nMndj+65fn3pBV3GM0oFv4oG5yKXsfzpBQatDSR5tVxPh/1AXxabxkUAyViN
91M+n86ZYzOwjL67RFHuA01SplUhSFxiFN7MKEIhOcZotkc9jm6b8Mq/PL2852dF90vPnIUBQxn0
u7xsEZzyv90acuYsijxBdW+RyCQhmpVzXbhV2QNv8gwMOPFLVxreS+YF3AEf2IlMnHF97lFJTrXD
k2AOaaJYi+7cMnemL0LjLn2qS2kDbYIFcjBtQ3ZOkGzeLbPtOv+DmDdl1YI7Vo6dXBVGzl37spK5
ozLAZuCBoKI23TF8nAKfTXGc4c9XNIRLNHl9wVp11yMgphtNSyiLCHLNq1RDiicWATG/1/BJn1o7
a+ZD0f9LYkYtBJ62sFQXrzRsQ8wLc5Jr+N3WO4/Hjt17jDt2z8623gRsB5p/dyVTaYs045l+QBH0
id5hxdpnZv8crAadpa7STQ3HKBz3xKmXoxzkILGR2KS5cOiZvUrSLUDGAhgu3ZRsHFAzw+Ypzw3d
ukjRHxKEuHQQRehg01J7OvNuTOQWPZzfq/ThhSqYWkISmcLO7Ao0jMo/rGNkghWrnss5r/VPjIpL
ykl0jASyw/5HFD674s5SS2IDswrsxRW19Zi8gtd6jMUjZpoerc3nrfa8KA5PyyPYraMG21tI2EzV
171joo2JHRoVd2YiUE5XIQPvUrhHsLaKHjE9PuO+kdeaE7sJGOqJtgcbs3HywGt9CpaDb45wdxDV
excys28NOJPp3ZvzoFNZoglaQRd+YGR2sl64J3sTl/YxbjUv9pgPjeef7HMvkVObp2lo7dBf6Kb/
IZcHLmlIrW+6wHKy7jb8wvosHo5g3ovhi0/H2EN30v/jxyQEWYxHA3LlwsflPaws3QsbgucWmyo2
a6Dsoq/aJFTJKww+lgk4aqtCWTFxtGRwHSjeETHOlUpbENohH8mNokhqoYKvyThhW4lPc4aM7i7/
vARsbjopS0xZ49oCYFy35IQWSHrCcvSnqi8uNoFgI9NNIF0gDADhPWzx2sezRUZWmtoWaj7NbEK4
KEHJJXm4JVy5VyqSkvNiHJxjCwdrhDC7cBpkSBLL1SCSxDiEkkOGV36e0CwaVR/WLTyI0+SGu3D5
bqPclsf03D+xeACd7YAPc7pb/QpmqUEq9o0ySpDRl3otmhjVsJwDpYCT7ksWUku4HC2Vg+a+jfCr
O5krsgOK2gnmTFry++kbeorFqJtk4tDWKL0arRMEICJ9pJu1+ijIG1i9EUsaWptwIqIsSdog8GEu
2dc9M6inkarFgu3eRlOu2AUbsCPKeErk+Z2vjl97qG6SafHxcyW1OvMK9UbSd8g7kpJovkWlg0cI
Ln3f0ANXQGwFZYMqJqWvvEsvp7a9WRhB2T/CB5uoxUzFHlgV4l9YVEejMx2oyUP4nT7yi/d0Fkde
7oQwFfRhlqeh16vOPATn2uOqASNEGEnhxI/ISBgMUVKH09Xh5FLT3JbkgCHtaYDe8rKw12RZTo9G
NTAgKoni+cLu2csu6Gg2w7x9oO8yKTtjrjVPNEfzrbviOrSdlnvRpSb/nTMa79LwnhsF/awCnvYe
cze0+29USsTSChGjiyRYFUPLbJ6nunaBl+rFMHjonqox/sIzGhT9MdT4wclRJ6uC2p0zbr8y/hKk
ZGpsHBEm1CerfbeklgcKJdljs1Tg8tmxMPfxxDfDvBdRCnec9qwwLJJXVtIiKMWuYbmcSjVa27sr
WI1OVFi4M5ZHlWudeeLFlwwraUP2mdsqbFu4kARfXy8ZtPaG4Y5iECiAVhagNRVUpdPbgCmUJrRP
jjyefYFuHsyWumYx9si346TqynJGBczo7TFPIzfVAX4OUVYNGnyqKjYMIz3npKJfdSWUJOIGv0da
W9gvDYrKfhW9bH41Bsexhrsw7gbB304pmbuceWYwIlbbLmLRNTpQvNFlCDqmIqC9xK1yTEQItALu
ohs5q8NZl6uHBijySpUlCjhocqVXvnlpa/cH2H4v5fsIBH7S+f54uPDpnckMMoPqUOmeFlTjGHaz
lXOmzRdBMZK4cO31BKZzH3dD3Dog0ZUxJOIwkXWUN5jqojiQk8N0fWEWqtmo7FPk6yFbIzd5/05B
4dpKcAfC+B0uTSfmwwl/ufsqL42HhHkSLO6DwJ6OmllwKAomrF+LwmmoXbOBrouPzn8w3zhu8Smr
DSToSkORWpTPHriIt6S19GH2CFNfDW8iVlIpw+4Fm0mJzT6eX9Kqj1z/NHFTMLSFVIdLAHixbJOx
F3aZC/V4yziQxeSYJTeVvmreT8V66oaGPjXnX/ckCESG1308LWZnEZ1tsdDXEXsDh5qjg+dFA4ua
5wExBZjwYo1SXIc8lNUHJywr0Bl8L39woGOnTCCAQcwEBHlZwBwQUJniRe4pzCnhZC2VSYJRmp0k
jk31bvDwDI8gSCnXLIyBiw6xNHlIe11qjN3DP1/MH0cfszM6maostCLNBUwSwkhWl2RtpCvBMwrV
d++LzHt2AAO28hX+vcGYWzdzERYpmlu1YYdF1zDW/T3n0q3x8ZnolO1pcnee8OHfoP5TUSX1WNq4
seYT9ozMZqz+1bh8iaqAmsZWhxZqPFz8Y9qY9xpCWMZdji3Nrj9k0p8JawMXiFGJl8UTUxmIu+rb
QVQKurb+SfgTJVJJYigYSskzP70Td7auOC0DXhYVMVeYUUY36gYSmH29SrlTrYfbuwU0kg8KU0uP
FbWNpasaQn0ndVuzHk+eCWv/wKBjy7ycEyFn/jC3UP6zPGUYA9yb/6VhcIFBOC6siTRpyt2Re1Gv
jgAa1gdx6Qcn+kCUe/C8IfzwR1zDTrcBH5S6bzCCcXrKlMm0eu2RPlci/YqHn3HCNHPgAYIA+0Hk
8Yo1BUhumgDYnu3bKu8bj72SLlkR6evtriAqTpXrM5nWFdqmX0hjTOLLRjS5YU5YTNfdQkg3HqmG
VxlRwk6OUD7wfbvnEYDoRp7Vf+JWffAACLX9XT2Sid1G9e8cQtr+KCQubfEv5GyBtPdb/popEmc9
dafZrsUIHDxqW0eHr3QyZpSiqynmTYy2592FZlJ/Sy9/tvtvCptZObG3Kw3TYyvXQx2aPFVQrBUh
LGIlv1DUE0OLjZhQ4UIofAB/2yfbO6ikJUkA6UT9H48QcM+zAf+98kyg35LW/+wV4Mp4iBWEseuY
4o00hx4K0Xpo5U7+0oI64NJvqr01tZNB9x4bbp/RA9B5MGG19a6KvSeEg8mQkPlZXX+qB/laxHaK
+8KgRtBxrHl/Uw7j9hnF9qZOdaWx3gqgLCQ7NYGVMLeiTiRvgyrh0zCNI8XSY7mbBfe3I2GVDqaf
63a8w6ajtjfhcjTUk//ZPGSvyEiv5T2KU3txGSV9BRLIFNYjY5kxt8X82tNEWT4g0jJfiUVFxOKo
k4mhbqV4nzeJ37r1935I2CFJxGdj5jzco48ssokq32FELaEI4d7xQaauHPqvxEN4YLdjiRUtn9hK
T1eh989xkOPdVeRrzbi/EEEoF4J8WxcEJ0uxqTqdgZ5gr/zQRe5hF6LNSv2D6Gov7UYAI3RzpHkR
RQa41d0PACuOc1tVRVJF4WcJ38YPRtAeeFe0N1RAwEWKNrvCAYaDd1RM2cO+vBZZZNgFfdaRhbOy
i0UOem/ll4eEKo7zw0/w5+6bQ073qx82aMO86BebqJmZ9oPZqifp4Kbd28jA31V6bSSep1jKZbjn
GXnQPn/83AtKFhnQk/TRELBULNvBUNxtJvV1iUqgSlqfk0w/gPHG2SBCiHCd+V/oC7doCT45nLUd
xSel/J5gYfpXtvWu4am4i3PeYOhKdAdEjsYCn57RPIQ3KfGOXdw2Ky5kmhwSrF/9AKP1O9ycAFKB
//aJW1FjybMa4OJaAxPH3oLtB7M7SFfcEjqRlcyVLGCudVUkZg7y/jivkVXhC6aXp0wkkXzMDI0H
+I+HuD/v23ZZdlMc+KKbFe7qX/YEP1vbfNZ01znuXV8+C4IwBh9ZPJEkkThOG97ZXtKjRtHx6xL1
H+uPtS4sz9v3r5jx2rXj2R7pV3mKmhuED8UfLXrhIelCFBof/3aR85OhHeFsHo0K144CFYfNzuXS
VwknL4tO4d9s4BsIHWvFbkKrAHi7XHFp81NURNKJKgkpxyOJLC184EgGaBBOYsbwpsU0+S1CPYDu
Fa4Z/RTYSyqJMw9hRG4O7059Kkm8Djpb/ERh9ap3db3RvNS59Rfe8rDMyeXWns2mT6hx6fO+2dkt
34taZPDTHgt2ZPSG19m4cxDr87ZurYYDtAurPv0y/8F2t3uRrvNBK+T8QOPC/rd66h+sGueFIQeX
JGbOy34cxQFp3qfkc0CcOn8zRMBi+an3DR2Lao7vRU+ZfjmU3V55lyHLnH4DtxaKnRH5vF6nBVgD
OMX2MyMHIE41p93DNwS/nhtBMxeevKalScfJH2eUNn1qaJaIScMDUD1PheITt5ifdZPNHzZIU8EO
6xIWmQRerJ6K6+1G7Joc6c1aIFSvJDsIjyMPBMvHHl2pB8Q3Stro/6P85vBBl53qjsfI8vUgK71y
xYSkdrIwNvmpLHKHo6uGi55d5MPmqMBAV7Tt/2czbpIyf8EvtO7OxyQhI+nuXlTSdN6mQ9Z7Acdn
PAdKZ1wsG0nFkO6Ot8S06wTmFMXj5lt4cvCitM3DuzUTMvrmr4DojVv3oVluy52KVrDxc2a7zIqc
YPevO49oL3IuzVBIQo0NQHJQ/YtGr4A4FXSingQmL14RsVoWz0XYLdtxjD9ciPqUgkw9Rd9go/vY
C98d0MmOxTaO48Sl+iqin7SPtOiLojguW6rTcPdPSGMy7AaQofr8TGhE/wabX4wMgyn6Bxqg508x
lIaBYW8t7kAj5gfFVoXhvvQa5AJRh1FfG4AMH/pcNudLNV/mGdcoNtz7ZWMBvUNwx7HYjU9nnFnT
fNrxMDNW5/tUxKw2Cb2JbfyjHedeP1q/Ey+J9g7rYgMgY9g9yXIcbdElJRDUvlU1zqjo3k3f9Xt2
EXZmNvl9dBZcl3pFAw6OuFPyMLnsuaE/9AMfOxLqy4NNIhSssdjAFHw8962YOdSDAEDNoGXJ+GEl
cMg8SFyRkLI9dHe71z3b2tqB4Pr3g870vaFIIkfLpVaxmyPxRHDjzuJzAUPCgSGs8umW4BSabEe8
orNgj/46KBOvrwQeRu9S4bB2I9AMJj80wqA3cu0J6qLcKKz9srFTMaZG3AofNMEFVfPyFn+1HSgA
1Bcdenpyg4St5U8rQ7UbwthKyI8crolW+w9g+9QgRBjDAsflalsR++TrtgiOiH47+YEMOzOceNDY
vKdHO7vHfRvlaDTApA2swuV4pxTYaz1EHojQ0wzSn/+zrM+EXCOYJ28kH48lC317Z9ZYL9/3V4fH
5Qal+1ZkutviPudX+QCX8HC6leYcv+DpASinbKGGDMa5ZzH6ImfEurVjXHGXkpswoH7CtkGp+gW+
dcAP6gRA6MQJB0VPyjGAAVp0zM54jvciRv+4c1I7bxpBdfElu62vw0t2tFd+w8AiPIWP4KcnxQWF
fOPaBsy9IxBTbFhFMqWtpStV/Ts2cZ8OgoXkhOJNP2/iehBC9IDC76Kn3GWDThJZO7wQeLUkw2hZ
VRiA5BRRaF98rEdc8LhGd2ms8eoUJ301J7IoKLUJrCFOCrOO3J0J7KvWUB402mBe7E9z81CsPt8g
11JcM7FB0lel+89cZ6m6wjjbaT03m2/ow6PFeWQ2CeCTwE5yaZBFbR78cmsu4MF2IBciHI2dNoc9
1hxxiTUmF8ADG6hIn6yX0xpLwmclhSNaQ2I+oYckzeMljT0h9SOIBcaN/6mJ7pI4R2eXyZfjs2T4
ici2hIYNvn9IJ/gv3npV7dozO2JoXCU4qbu5HNjgJFpYci0mf/SCnmQClmud5oPb+J7ib+3bYkIv
ZcF/+tjAkDsLvWrIqHdBJh92ayoAEFhtzvoA63icSrPp2zjY1ETHt6CwW2twfFJOUyAw13cHxcgo
zmZy5xYaSZ9CQKmv9PxbtJhaQLwTTxObkN1zQTuIirgm9Ntgnsgr7Cv1U+FMyFnCCFnfGjSt5NQi
ash8Q4qyuk5SBHkwK4D96j6h/e5xfeFVqzGKfxABJdS5MO2raFXlYrEsPdu0IennuEM8OdAdGAQL
aK5zWvxpU/jVYwscyvF3nzqgw2X/ZtpEFjhvu/XkwhLNUs6cicPJZL8/yEgtFh/NIwAhl35BCfsJ
dgBmjGCOCdhG/cSYIl55ROUEWA90fMSXpNk96tY853eHLOizmXwcBUZhPvjqDz90mypG0DfE8V+m
siPpHMC5O6gz8QK3CcSePvXEdDkqMEc0bxoa1hfbE8M378GVxleb6zSfxRESuef20bXmNGpwKQx9
65gATQQODR47myWJNWUUoSyGCHRVUzRh/Jbd1htASzZh59OL0eFq95iCX/PxQDQHXXWlASrl+fWH
HyYE+SSE4tkdy5fkCaNTzwJXU2dwNhQw8E1UGzWPe7NUIuX0ALAfLkvu8EhhpI0He5U/OQHwZ5t5
hcR9840c53N2kKyDeKI9QHcLQUd3s9X5cq+m7mZNfbfGe6sfg3oAARaui3it0E6WSqlmu6WB8HJD
BALGcgw9OTVxEsqv8wPlQnGXnl5pLeRzx4puiNY8SPfHPBNjSsEYuJP89K9MpofGCb4QrW440xcG
M+8aos+QRHlJwkQ5Udxak6B9A9bhfqIVveX54ZOt38f3K6Dc7rpL/GTzL3YJeYWStCYhFHZDUtho
LBivYBBg2obmWnjS5r0yJfBzc2N4WEaqhj5jLZ5TlohGHcKzie9EWN7AQ5XjPxnM9lNps/Axv01v
eBB2G3Abqm91CG85g1TQB9R1JD8yUnP6xXLiubk6S1S1wZ2kxj7vaTLyJvRW3MnUubmevFfm79vF
cp+Bj2KsYLHKts5triv+0shyqiXtN3E/Va4kZT0hBx/cqkecYoK9SEuU2u4xBGuqJfsvhGYaBVe5
v83LpTBFBKyohnp5lHfPkRtgcjbkPnUb8U9TvxWqVXDZEyV39Qq4vnMq4sK9Y8jlsW9qap4XnDkl
GAdUFJXh/BfSSu0A1MjcAROz/WEP7rdUfLxqrhixbklt+eiWvva8Nj4SVrLAdb/Bnrmg7uR5MAuq
vBH1qwfTH4sjpk/OW1RSArx76HvZOP4IBwwFTI5+I/kakeZApt1ZqYY13VTInXMgUZPvNTkZAdLz
HJBIwedOChT0XCuhE0tLao3cpNN0uj7Dr739BnwwP6GHiwRR5R1gxhjQMQdGGme/xenCGjQFRYvM
cElCXESaxqilRHKMQzw+7AMgGMlZ/4Hr2d19MzUibp5lQsEOv0YRfAXJ81RcIYB9a2wFm9LPqwPy
kRr24BOJol0giyxR8Kao/OsAIx4N9lpnDvV5ZNvC2RFgbeks4ls0nYcmx4IkH1DzJQjgdZ9IiVTW
PFAmPseAhGfJ/H7kFWlsyMvDrvLiUjLpvtqwVe8EyEyMFrDRJvkCK85d2J+BNSunSLCrD6+i6PxJ
jz1SH4lQS8h0Q480Eap1l2hKQhskLJDgDn3zurokBpL8ZRcUkbBQISSBr285mZIOkOU+nzUKXhQI
wNxu8hqxwRtWfCgqQSSEzCiGC/d3QJzL4deRlR2OTRWgZpylHhImZyTFCYDSQN1viNJ3fH121gEw
SgNnixDB6hpwii66TM+vxHH8ZfKDZzhlH2BPUhnt1CCbz9WH3H9HJYTD3/PLkpm8lqFbebqeAJ4O
58+/DYToSSbDrTbBmljcDB5uRoF/qQroTCjY9GBKVWzrT1G2CsA/AY5/K9JHohxvTzkBN1jiMyBQ
QdHuUyBQOURevYC506MzfP5n3YJBOyNPbTE6aWnSw3S/cAXcsJDFEhEYq95Lczz2X7Tq7W8720p0
kZHhiiU+tpEv32KBdEtho+6XYbMdL5tPrHX+CI4rQpUEUbJk4DWk/2pV36TX6ZAqja9LUi1Y4sxC
J9N0lXLqdxPlu8oNUa70Vv4NLAUnY0sOcye2bTRR3hJXCb8lbQE8rTynIIuByLiI43tp0l2LMJMy
dFvBtoHGdnmL4fxKvLArzknqaJCtXbmZU2i0usDJI+yUJXEwY25uhTYfwEmaysrnfuDr1HjBp+y2
1MV1aLqcQ+yaXf035UPzQRZys/Z5ucfqvnF9Bi/3BrsBtix1hNZovA0SapXhuNni0eUBxoBfkkhy
b590uk7mjGTpi0JHWjON2VlD4a152zzWzmANeSiXi+ZOeZpjCWN0dV1YiT1UZmNeOtJQYmpTi2Uo
y5Axd656nOv9FSDwKeMVs7ACd+PciwtGV3DKKHmiizW+d4KghZzdgXjsaN70xGgnP+wjy/X0rqCk
n/1qGOJlCdK5QXj7Hvvk0O7TvDJP0mHIPSizBLWewtkXYssN00x1WVg1zRAGmgLFQw+8YcrKWMt6
zk8IkSgSAWGfUtSpgS8fM/zkM3+akpO3Ss3k1v42DaG4sbL4kPRhN/t7M2bANPbAPtlBBCchgRes
1kyrIgj/tJLot87O3Esrvot0xoMKL9UMRTo9Vdn/UtqhLVsJ61E8L01bX301/Z9zd81KWA+SjzLA
MOXg8NFFaml5bD6+i/Xch0p1DfEOF0S6VqNsCQLURq7I+9aha+KaMtGtLemhOgPqhty5MOJDjNcT
otp83+oPC0rPRvM2Awl2BCi5CvvuEASrkq8ojH/xIqAor+8VBBiPa8vYERH30V0IC46Gv3gDoiyf
rTBOwsu0WEhGzZfLm1SeNOKUGxxGzs0EohM/zC4obWRI5FrqmPRvrzlrgCG+V499kZhbKICtfNqm
kf7ZCoucAP06bDBZlAaWyzl99RkyicLD81PjMwtrVFoFps+Wr7TIdmsSp8rbhG74h+GFNLskL13F
Iob2DMja0M4W+RqRU6aEvz8/z9ZhW3EKayiAZIcPa9wya0n+mdj/YFb8ljcn6Tdtotfn1qCr3JwZ
puldT8cOT74G28zzwEVaTTgO8CboOIA9IxOpjxuczUDgq5W2sJzrB68iDQSziBvvNVVuVUHj0pVI
b3XbA6dFZMRzDdCpk7GQ8nsymHWQ0ahVNquDAGorHZQizBI+aTxWb43gvYs4G/BTGajmj1hVVSlj
4TSoTqUJo5ol1w3q0UwI1PkbiV0t1+jxKCC/Ag+AaOEDvm5alvFFcaYWfNVsGBfT5J0l09fJ2kjV
Zeaujpr2peIcquaqUDiBxZABJd/my4PfMsqQs1Kctdn/+hUFYL6shZU3V0DAsa6uK9Zbzi/TOcu+
SESUmx0efzTp5pmgC82oNROvb8JUhvgSQaY/h+Fi9+gj3p60cRKFHYCV0uoCkswsvf+860zw8U8Y
0v8mWlSkElbW0jHg0KOV7KEpKUfjueZIvwyT/DsMHtyQiaeDDu0FmEqy2GWbB+OC9foy1lB4/YWZ
IhIVSIG+doHYnOKVTHE3p4US/fp2xJIqO1aV1YFXUtJkboKPHhzjG6v5olO4rh+SrfuFFmWp1M7/
48RmzUDVWl9fbe2oxDiGmk/DfR2Juic0TpjT2/UAgmhT7jOVGM4guGV0RamkexYeKN8/q+167ph6
hgaCwoh8pHunTOVwlUFApSp7Upo5iLo9myl/u4VJPTgi/12HTUr4SZk++ourvYUJWUZ3nwcQnRLp
ze6rZygYjKZKg13hancK36SGKEQ/3uGteMpXwHi0R8vrcGw3oumNywAPl2cf7lbxW1cDs9HYQMJn
PI7DthsYIa+Eq+3UJslBn/67XhqQzMGLStIbhG6IBNF92qulentOEFWQOKtyDTDQ2TDTwAWWKYoA
+ktp+dKZIbUQkqssaxrMMd+NQhWNRnVBeOaqfcLa+rkooC4o1YTRBOXbEN7Fn1FuM2eqoOoWx4zd
AiIAwXzNkd8WTtif+Agt+7s9LDEMCo9tWa5HuzdZqgqtQKkUyNyAu8v1sAdYS6s6Ow+i8EjnG7rc
rULS7Mc1qYTbPf9ZH6GEfzEh49invwyJxnQB5bmerxKoyb5FWDKZSOiI/HuI1FA3jOj30FNUGeh9
ooXAPzcreaO1+y85i/e4gNHu/xdtAJXAr673xlxyuoy1gctlUlsldrYTqu02Vnn+ZFWmZNLXHz53
AH8kRZQIRqi/U5bsvDKghagNDr8fx33ng9YLrRgaXSFOWZtGYeg8KQqm58zIx4buOwiGeR31qIkw
iic+5FZbmim4EtRulTdtghaKhqwCE8vSHXhwJ8XQ20lU1It+76xBVDdAYGk9Shzy+/lkFWIlbLw7
uf/oxSh9TSqS3Vu/L5LH3YOCJqMQVpN9LP0UG31TMf4pZ/AmzqxdgtmBWty0CowLRoVHv+AHgj/u
oysmp5houl3CNQi3Gp0SpFWeth2GuCq7/q2HtNE9AoopD37LIM8tthwvUAMdp/++/YRzx6+BT3Cb
cWdiJFhXRa4wXuuI43AXr4dmL0M5I6EJZPSeAFVPl6pckT6n8pllTqOTe6J31QFCfiBVZMXWzg+7
Aw7/W1SypQIBprGC6dOnNLSrl771F0wI2sjjCHLayZAxVMugoapmofTCHGVFHsPz0KWXFTx9p1YD
lzoCMfkWQAVRjZiihpu+dCQXtZGLAUvnGaeCiAgqJmfl4COc2BOsphK/lh9TRPWcQlqxed/qKmxw
lKoQihEb9wQMGu8qmN3e0ajK7WDmg0bVTyvoerORHAbxy8d0LCa/6KupvcNw0G7mMz4bvYBSxyGr
fWSFpUKKHBkl9Nm3ruV60ndHS6iwFfAAvp2c/b0sSZpMAdAVpk0ibKghYftrBiHfaEHFPfhw9BR9
h8i0dN8F+a+dcY9cIfam2Unr/rRUG6b3UKiX9vF4lO09KivVddNB07wugStZc9Qwk/Lr/iTci5A/
CJlIGWuD1n3S88IVbGc4R5+Nih3X9a0/oo7G4FBsgfZf82ZFvZImyxJAz442SM5sybqbqac2aIAC
AOkClH/3ytgXWGKSujWWgH1M4sw7A+h+OEx9k4ZXdFBmpFY2qqWU1fNEKIa9lB1pgyyingzR5eZa
2gKX2wtLcuhiNZMOpQ6/XhhSvL1TDRVVBPhL1FcIxyO3aZckoJBr5WpgeIfu9oPc7c1fqR3BiZiO
rUUS3Azjv+1Mdl0y4vKAxrrcYfdzmqPUsQ2EkQlBNNd1oDiSly2o3p2fURSEzVynUeQ8z0o2ClZ2
Ri08YkujjrieyVPgqp2xf+7YfdJOUEfviS7r+w9sT1VD1CQ+uqSwkwo8JwqdRLGRlyybxVBCbZ5g
qnwKSPT/5bM0Su/QPgvPwUqY8swOAkoDNyMfNbbAFh279WscuMOQ4OQepv7a5iw4J8YeRrSScJEW
S4ofofJLxLGOBitWXhKLTu+pkSmJZEw7vX9vb4ICQOjsC65lB6jrDxsyE6ferIDYeH1QoUhMgjKL
rEpfQ7ME5rk+gfXRx1WuvRThBCFsBa8EIfeHggGOwktv9ca8GDqBZ+Us/rX/uKs9zpDD0lkN0p6m
pIfI5a4zIwoXuTwLb0dNujocmags1a7QiOMxohNYcN6TFCKE4Vj7vTUeeTrX2eKK7+s2RqcBByeY
U1SbsiPgMUYbFmRdKbaqByW30eiR2GQWKglyixs5Sq8hxspapRfrMd0eM2Wuwek0f/C+dPpLLKWl
4SqyB5zf84a/+qlCY2ETHfRX2YZVF2otikS+rJL0yVDkKJY1MWOFtuygZsDTdxp/YW4Xsb1AJ+3g
4ZzR2PQtdv+rpqbUw3DDSmScNwANA+MXi7qt7NxwMbBRvGja/FbWmba+Jj67FJWKHxXMj2RV1oH7
tsdWTt+q29aD+eFC+HWYgSg9OdNOmtaATVeOwkb3EHPzWG7Vce28NqoaLOeaPOjFtDPb3UpIPBEE
5MDaJt42qcrQUJWbqGhkQm4xn0uCyE+JDzxuZTYzDMKM17Gjm2In88mmhMc/RUEpSk1bUiT+VYZX
Pr05j+kHYfzfcVVNuoukXE1DfBo/c/axoGh5Prk2LY7QhWBuFtrRdGEqTwhkWqe199bB+OwVFIS5
Z7UUYp0kEOG2yecDTBXYYpIblScw4To83Lgm/ZeoefDcDXIVOECDi2w9FThjaekix1oB9p2nS+sv
oLBj+xFdL62kC10xc60/8TWv9El69nfMhrR6bXxuNfZxr8DS7inOs+PmUhoC8QhGpVRMyaROlwCr
HfMvnx30DmkBEU5aEaNP+WAvoTQ9VXImZEGF7UfHz+biQhkBoQNteVfDXZn/vpVXWLXLOhKvFFbA
EZnN3pULdPXh0PYLbh05odFLmBcy8B/kBPw2wUXx/CoaoBYxNTS9bY5lgUFq35xJGEdzWgqH8/pi
StqVg872CuDaw0ZXxtrcmAthhJhKeHH8xYNgmEjA7+NyQcfmVu3eZaPEpU8g0vaPq/esJno3eqyf
VtXUU2JAPQRMgF004bo2WV9nq/YxCJt2Wt3ftU3ZB13ta3HyzGV/JIt8dRPRku48wj1YHvlBBW/v
iCnZbrWt5U20tAvBmHugj4yFvi81ctAjrJv5IkZ6P45l80T22qDxngU5uKwehTASHRID0+u9VIit
3f/ImNsV6JHbsxIoZb7Q7/FvEe6nsIidJA27UepddWtWSeDI473gxAHs5jO2bPC+AGuY41YbyHnB
gvylGiU8fRrhCSxE2Eq5AX4XcT/12Od0M60MDSBIr0P5/NMSuyCcJVaLEFN73mDqxMsIMaoPGK5u
QSDRZf8NTFcc7BiPgD6uA7hqUCrgN/tjDLDGBhAL/PuD9+jplP+B0qhWqz3IHyfAYtU8CXuFIefq
RzG8HCRBLFxO367ZHGSSuaQto8y50WqD2g4mHs1AvSVo+fmnOMI9iClEn4f9Dmok76X9BfBJTkYf
FncM5wyatoe2h1lvE64GFcicUBG1DZMEkwEMl43XSIhdfCuJTnfUPqnQzRP80OnXFxZEihIMYcxU
6TYZqiW4osRIGdelcyZYeHKPbEfcRgAAUr4mpvGxh0psCLRb1bc/uDh1URnpijVq7kap99ZTHSn3
B7bj7PCol2lGEVFd94exG9ML0uOHFPUZKML8r/xS2DqmnWzwXi1pFuV6HxrbApNociy6roOHp9KW
X5Z6/PsfYZRgLFxCvs5GAIaZrATYQxHpXRsYc8OfXS8zuAd4CXQS6CINrAkhsYibCYKDo1jBAO4I
S3vfFIcK+/UGpgW7CX5qrNkb99qJKRTD7nJajJE1as7XA54MUTBTkE3CThN6rNXUHeYpFIXkqQMB
eRNw8Oy8YoSC7O5TzCuSt2rAMfSFSQ/vP9+f3QRVIsEySDElRGNiLDixaJMBvYyUe/HGzs0GIiuj
aEkYrB9t0gp4J+gkQXDyadj21a5TtS+CgZNzjmFvP6/N6uU+gYhuRf7XJfN8hVSAeDf+MN/DyNPx
d9Cpz9tvs53vy4JtLAagMpWAoBx18xI/682pub23dso0j9ksShSN6NqnXkN5Gad4B4lCu6uQsYjO
h9XW5C7kMyaW2WOx8fACPkp3VO3baIouvGARr5Azq8iiJbVDFo7Ug23Iv2AlPYMEozEqs4Qw0olh
iMsoEQcC++mAOwiVaqFjsFNlFVmRKCstJR3MlrrFeaUfRO9mbF01BjVratGDTTKZDVfLciTbtasi
f2CJp8eNG3gEw0JI5qma7KnPykL01C3JimDpHvLAETDckY5wGHSlNKvnqwhvkhrRWRGj3YCXfrQ7
ITN4zc7zvdK7qKlBbkIPSUlalarglFERTERNg59ArOr4awxY2gz+f5Ye/U8EyhIYgtufs5FheUxn
0Y7mdhftJerJX+fXYTzfnDQqVjCIZ4Q37Cp+58T0/r0ExFC+MSRQGXMcsKI0RXyr9fgd2DTyhAI9
g2P7bUmsmybh85aQPEoJ9y89RmwEXklFDV6oIy9yHNLbJGHSFGc+OfZSG8cBCxKLOM+z+cGnAG8F
eWUgXTeOuLX0qieHTnrdhNujk3De/Og0z1T+C+rjMBwtcbI35nt8qDmxvMiLqVbdhnqYrPD+sMdW
B/jB7XdmvQscR1V30Q+LsigiFo8Z/hTUzc9Zx6tw1TRjfug0W9iIjEELpLpG4B7njeydz7ymib/l
rKiRcIzeMiHxSYxeyK3ypPJ/HhbwcbDKfxPzH3TC9f2k+8g1QelDytF1Ao8QfajizUMq0+LQyUql
sisYYo5HmtfldGIN/cHfSL/Ef7pLc/HrTDnGalWIv2qVb5ALcPeNKzIRzTpg8C7dfKnh1yr6vOFM
szHnDsq8/M4Wum5uSl9A4s5bgVC83QK+0neW7pUYyNiHsxGUo5M4k1uQ7b1sKpGRnEKdvgLZPRns
vFa9mXZ4NTI1ikZje4HaV6KkBV1PVQyY2AM9ErkTdal9/+ZDO5drjWGD3ZDtz5B07s+ds2Hg97On
73w4COtbxZ5hRT6EwgVXnUvcqADr0I65XmeEUcXHbt4K1dlIzu3qk6RNsyoKZ9Uk+cUubW7s1DHc
YmNKnvt4iOM4/VO+SgIREeBgGL2GoY5xumeQJb2syp2kMwjD+U3L0SqqLbKDu/BHDjDxQrJlNEyl
KUUkV1XHshy34St56e9y9nAQhRo3hm5pUWEn21w8mIkbA3rX2fwkq1KMA2H+8PCUfPXdnLfD8PIY
Edivbm4TWuLZXh5mmHBWb071gPRfpaJxwk6wnkgFDcTAsDA6VFV690y+6wo1vxFDMuaCkHOyHtqa
rDU6WbAL/b+zoULsVzoHTDJyTHRrGBlN+nuwhx8XkfK4aUZxuQ3BJAK+ciaJ9iODFdMTziIgEpfn
zm6gl0roatXK5iAbqQxugGyINcRwyMIgBRKG3cqhwtnqXXyj5WVRAGYItdad7B+7OqH/RilU6ftq
rGnw5rMw00c1qEuY9D/3/LVI99n6tlAv/8s1IQ182Fi/HHqE7UpVHUiauoCVfanWMDrauQ76rL2S
RARWdydow+hTFT1TKfMw6gbOscDN4CGSyONK812JHdOO+I5UXzWJivBIG5T9Bi6Ib4O/SlkRarQA
/83fqXLYAzR9K8n4P9bxBaI6ISNeUk0jNhTKxtt1rT0crb7caRWYvbhnXGfz/RouEEbtfAB6X5Xv
bfCiqzUg5r4fwKSIPXeH3kmYWdp25Euv5NABi4cTHnai/raoZ2/3AY3dnIIBeZ/n/IXkG1Z62m9g
VDrtsQsFEOnCYtVikCQ17M5o5wfQODh5ywrTXJIs2XTsoF6hM+jU3LuIFOwk0uj46MDUE5lIeLa6
+Ho024IrMyztmQt6WC60Z5fOUQbKe7QHCfLy+wa0TLo3eA+LnsqMF8MwWPEbdxSdzGuujJDtyKoq
S41dPXi+fo8RCvDGAWG+6Pp7n+JVPtISjVKvQlCDlLypNYSFvqjoQ6XtEH1ixSXmbUt9QpPvkqgE
Q5LpMB+FfXnyth0wsYao58k1ETZZElLFtGNV8WEaZdZMhf9RigPr0FHoxJKCsjowt3TgdYme/FSi
+CZutr4X4IzOBEt7wsRQKRbObzj0r9wi/0SPEx0Un0P2DiPFs/gmLGNF9JlFpQ/SmcyCrq7eDZYA
PKsHO19cacLiRsXY+0G8v47UnsTTmMZ87iDK2ggMd998wSt3OAiw/lxiAHMzTYJAgA3cbPrF51hM
V5NZc09YMDK1YqdZLWfxdi3GhHV9Dfu7/i8f3XlCQqnDACXzwFQL1D4nyelCeFsRl4Y0c0wy3BDy
82gy3v93W1c5gEpoPJyaWptNgHSYBy3blZI01ZuMl85S2guSbB/IccRvsud3Q6OX0UYPPQ67iqB+
+YnHawW2fZliLVfqQFsdk/F2iBbgWgByhDqf8YKrc2n4DBNuFRo9i8lue1N78zdmMzU4mQyo7YV7
HSUA9mi3P4IzE5uXkOZRzqbMwQGvmc91A+/BjLhpM1UQ4O9xiXQ3VIQbEQZQnYzBl/8uc4a3wHJk
norEAH/UbEhA8NC/x/Szwhxm0YvP7CVAJtpmXj/VMWw+MwTVXtedIjpsqmRg/OfigN5hNGCEJ4cN
/9dKmeXZVw4blA+C7dhhZ3oP2tOYmieKLNRTX6wOjrY+XzyrAEgPg+Yu0anzOnMyMidTsApWR5qe
t0TQ5XNbBAL8HQJWmpzVGqRKa4sYr6zG32nGGhIDxp8/3z5K7CA87bYZ9HRTQTL/7F6tJUHF3wak
paksQbm2dM/cURB/GyqgAm4dM65Q21cTt4Fi9sm3hxLVEtLnRkJSOeXL6liwNHX1JFNfdvybg4+3
9zKthsb2j5C9sERuTw87uyhvMr1dNCqnZ5E+X2hhbbRE1biVjta6FUmLq/NdKCJGZPMrljvmc6VX
cABDkptjKmiiEREiCtl+W5BTXqx0kG7otF96DjM1/NLt2qz5Eft3fXq9Z+lwrxOil9tSsntzG5su
jWagZwW5nX6q4dz1ck6frqklDjNSGOQ/VBaMh21cu7OB0tA/p5Q5AtZlVrnDTFjQy2VBckYii/+h
mJlVzG3v5uOQ/kCVpFuDnySGuOKUATZvPOikwxM5xNb9HASzyF+TyJnOTKnQ7+22573iK3aU7NlS
cu97RuZuU7vitZE2MF6NzweZoUSO2P7IMeBELWPLQGkDZBFcBfvufPMtaKFEa9skh0XPq0/6mMx2
zAlrtOfvFnhSx3fQMwvX6D8RNN3ZMpZWJUJt903KwcB+56gzOsQpFfPNty9MogumXHUViexAztBd
cGOH2ZfcLPoARdiSFjkrGCGCLzjm5GOKkghC175OHqmFzKDO8EHAokjhPC5W0kmG0b0AxgiEAjFW
yxUz+ZDrtmPNhXyphHlaU3r3RwoEV0BGjscjbHNS2N/XPpfo0Su8JTIMVuDGsMEj3sGJS0KjoqK0
/IKc3eN5tFJXRVKqCarMbYlIwm7BJxkd0lda5XynwYX5DsEB73hCni3QVfj3Cu2iyxdEJQCRkztH
Q/ttVMQvUJtGvjRteXdDm9LQctAgQHc9zwanHO0LtnX1YbRlLXaWX4W5pE/Y90rarupmox+xFskT
L+CtXxdIO1pM2XGuEVJKP/XouGoPsmjf7hHK8oRCLQYLqBH/SDgXRtr/GODECG//sU02uHz4r7uz
wmUNQIpS6CfMoZqA1mM8l8q3lRdSU5XjmGNcCI9Z1dAIrcmJmY+TCFsFU7FP5n1uzsOzK2BizuHW
8TXLlBzOVW67wW+WaQUHy9LCtoPA/NfXg38tyG4aSgXe7oWnAhs+NQPBDZq43kDOX9LPu90Kl3yh
lmQywNapo+3YVhxOCLUE+OdyVlSdSnRAUj2qXSHPYFtio81ox9LnuGCFdMYYtUGCm7Ka0K799RKx
hrDSjZyxJhPw6Trlzd3ZI8y/1Tmg3AClYoejM6yO2SKiEuBJxSKRLLEM+iC5RirZ6PuCsz7R+FMQ
5FGJY/ynoYYyAUN4UEC8cl54ZIgr3j5b1sK6ZiBIw2ldoNajWh0A1EnDD8eGC/QxzW/C6ngKTWE6
HJl3Q+oBzYJ5Cnrm+zsoRZm0WgiYMFDoNrbGNxdsUEMyVQQVh9bA3Pdp0gKTNdxZBcSnYEJNk1h9
X1zt5X7IZTjRvA0NPQHYEwDVv6iFxXAnOTa73KmaG3ZPaS6ua+S3glD53KOrd9xRnPYXABmN9tsu
VuWlSH1eC3wzSoJmYiolTPoL8dBf9NwTEOBqWn7Fkkji7dnE73Ks7j50ORWTzlK81Ptqi/qUPhY/
0BvInGebuosD96KTQMdyelMSGNxF/2qf7TU9X17nF5Kqi/q7PKvwSQQ+TP+Wn8Cl9BzJBSmTL2dy
uIJ0PtUrtyubrdhuCgZ67tUUbU0R9WSPjeMtFxbJHOl74TpnZ8cAUKtIOpfDJXoOxe7ey/ngLwJZ
nnURzurSt48IalcpXHt0hVFKimJJauqvwDRDUuJRzeohGLo9oDKZHZSl6+wSR0weOmCm3NWD+Ogc
RnVTdMhsFtI8fJyXn9fKG1SA7hws2irAHKbqi4A06gnsfIUUepQeOSgdNd5coISWXeFLOOXgMtd8
vrqkIioJXRcXiGqXu18vdZQB+R/eFdF4xmuWUCqERL7JuOgUrxBCTmmhmGoGB+1lAlcjE5K0nrtg
GwUVKyOALiI7E0iX9JgdsS+yrRheM6BicmKW/v31A+h+ZTjQJDGJ0l2tUUpf3lJ1Q9FB76Uf1PW2
32MkWkC8VsElJsH00hQlJAwaCMz+KEgaC9u+criUsAq5fsDGbF1RSbzhZbweK6oemaeE2W2xFYAf
8oMMOLSFxDaibEqprnEFHb/8VUJRe/XrUs5qStSCAkh9jZoL79IkZq84FIJ4agqe5Kukv/SFQaKV
DA2WxzgtMBbzHtSdzOtuQa28XCzJ8wPOLJCsZO71RMme4pB99VcVbdfIgbcreMo/xUlREftck0aN
Lhdiyx3BvfB+RZacpO3hWXQUTLFedIZJ5tV+v8rDt5kiiEMrIpKaVr5SgvadaxFsUB+DnwtpGX9x
8Q+VhYBmcG462+NVeGRukMHA7ZCTb+ClUfr8vS9PxMdayPDFyYfrTVvHSOdoKVAJisxkZT+Ap8bk
gqrAPF7A/DLWYKARL4JLOG0MJhRRRloE5G9I3srRvKqaJarrECJf2WqGcnf+SaYAmO7outvHi8J7
IfEaaQi4lS8h7AO9CfL5qL3jV+CbKVxPtPFWyvKjU9h7HWEwD0fhGCiIKXrt+eSzonrTHIQHdiw+
jtCTDS9Vhs0i0g83zxrNC4XEQh/fuldCMP4v1uOABgQBAbDP+xR8EYPi2EGyIffnXRX3qC6DAbvr
COr12aYC+1i2fMLqrxurPCb7rrKD76DwNoQysBjF/4PJBQOizyUZwD0ktvEwR1Rtu3F8pzL/JMEg
FfnZR9fMLPuseIKpY4u0CLEpOtODMEC8JegOAp6GJyymbKsNB5AM2sCBrn1F2oeOe8uF9pybTSk3
uxn4wYxhyLzhlfVo2dYxXLAiblx0ZEfe0l1/nE27bps06uSknRugqcWaID+BcwvzMPo9S0/CIQP7
9PLJmXg54PZyeoYamYJ0daZGBKICyDkCMWiriFV7IChU7dbA/39Y1hITXcO2O2zJN4JkjtnrhVLY
2vaFJijjIOc01cWvrAY6snfCqdoQsbCYB8TuQFvFDygouzeOUDrVolrIyHzr1wp2TGDQpNhXTPx2
A966jV7trDp1H6SuY4Y4XA3Ei+B17tTpu7V0NqRsjkCH+WPfzWuW4/+DqN46JVDNpZbKMYpLA3Cu
sOiNbFesKDT2VoKaszUPJeb9IivferQsBbWRpf+xzmyJao4q0B8Xtaf1vlpakAUhzWYlMx0KDLcd
2UMHCUVqDaYcoW6GhELXNUjKn2B5v7m+hltw+Fn4zljA1JF++TZ6u+sE/6K6/bKpAYS0POspmJY5
B4Mh5UXxi0bL1soPy4IRPZebzGgZ8X/O7GAE5p58EV50QUpcLxy3S5sMvDQVAv5xidwbVyztgqkZ
BJ87+G+US0D89j4pfCJQLca468YkAB698HY7HMAtS2bKLyc2UP4wBTG5+Zw4dp8AfFp9uSRkWc67
sHKzhoybCbWlzb7Xx6aU3n48/y30vevtQoz40dsILzDHJuHG1oLidGAV8EpXOyV7VeCbNpFiUfGB
noz5tnQjri9977LgqRXcuW6dNbWh3pnkQT95iZCOpWaxd0tYBgMxDaG5vj/ujoFz645n3Ojo2tGL
815RvIw/xNMChSEjdXJybjk3r1xTY5f8ZkvZ55XAnxGLo5E+6LsV3Fa0V8G/OQM5Wc0X8Xds0T03
+q014lZzrsHmGzuXsWchHyQG/lHVMZ7nviCMpeIhg2ERPKtmsSZohBb4mk0hW2GTox5V3/GoWbNN
cfm2AFvFCGKd96Dc8IlEa/lzHc9iKyRh/bH+bctZvDWirBiSnd/qLY0CvuylEw1VV172k+yuvXVY
hVpOTGa20/JObfBDXvXgeXhyqTP4ZPYjC3ECBM3enyuXaYhCIZUqme+RhKgpKvZssnuECJ7xDKSO
v/SA7tHhfklV0zf1jGP4HTRl2oE5t7tfH5RUYI3Vfe7m7wReKEvALPC9izg5BUWPDtLi8x07s6KB
3PGoG6bBFcYFD9PxjHydlEHhOmZLAHV9xmQZENXQmI/8KXQIIDreH1u4tIN0Ik+9d510yCVuHIHh
qB2FNw39R9AduV4VufQEadQnl8+Bwo30wHGZfyoDWh/lUHmoiCajormNisdgAK9j+Z/SpOYc0Hw8
ImGUZ9n+NXgyh4JEj0kl9iIJwpA29GyIJNj9ctnZkS1m0gzBJ60hGuh+tpQ6lFcuizLmZ3T8rvzX
+54ZbXqaZMxraR5UZ0Kke7+NR4TwQegAORNXgayFVWHVxaTDkyjkYR2H8ENy8McoVJS4F0qYgw15
Q/8OZIu6B5hIdfECth88YH9387T7zC7ZEpaQfY01u5totNayIHcoUwZ4FYlb8jsWq+IQKS5RpsZs
r2yWrLk87TFl3J1VmgbCggTl9/od8FYtklIFbA/LYfoPBKzqHSpdRs8OSN9r4RkIwkWC88J41laz
QbKAIxBXiYfd9ZUQXdTVI7kXutJ8IRNYDdnhgqTrSXJK6vnJYTLyBd9AY2/bIwvexzTZOqnnjScj
LimKTicInBhJKgZya99iBeyMNUOcP6Nm3HFPUBc1xF7MNeKtAcYyBllALHQVioOJG3gAb7gUyDPL
nQB3Wdy1utPCe4Xt19jN9RsxYxlhEGpI5oMRuQfycM8FMrH/T01wxdnQkIng2XruC1unkTFEqRv2
t8YatUNfs4GkvWBBnf0P1QKD5PGsOLUPC3IU1yh5Jw1UDq7kJJG5ZClf8E7WNADH0+jDDNicgGOx
8PWdtzDr2xwOE8aXzWXmPfVLdUlDTjK7+g/XDH9DJd33Ke1tYsMey43RWKaX7FmgOClfwyRIpLWV
+Q7WO/nrrtedu9rHL9JwtNGCNRC/vZq0F0UVSNy34wurljb8kZnjgqRrHOT55o0NfCijYfZrJIYE
kxTECjD3XbXZYLeOa0K3IEaIFgj69h/K8tSkLVYYM5T8OmlUOPHVaHmrd0ixgXs3ob5SDBGf3Nlq
NC/O+J/31svzcWlnwpvS9yxL+L4C37KkyzEkmZf5eZfNf/XsT8kReOApkUyb32UKHjqp+bhNpQW9
3/51XwkoPSFoL/hPvFDlvWsAizeURPDGe7/uloG5v/cN5P3qLdKl4Uz1N93bybhI8RrM2IcjGL//
Jsn48HWoxdVlkgH7sFRcOwlqYV0LTc2Nq72lPptSvvrQ8IdoZXQs2YLCYCdVubRSTDNpdbijSZIX
+FmuayrJpgSTe+FmdsQdiG8Tey6LD7P4eRJBpPuLgSxcNnvbqa6YjCJM6MWSzkXO6otXw9tgMa59
k5Hudm+cld7lmJdlPN2h2WTI0lythXbhWhBEeaXaagssC3ptQW0F8HUoJSMRoFBEx9/DbAaW2sHS
UQZ7secUu7IOGZjPSH/mFfp33mPtpMao3aKOj0Txx5uL6QBUBA2WN3cyfjN8LFN7e/yeC/RBxaA+
3Fl3G+B8BI2/TLQUsSjKIvTJcQC625ck8kszPpwT5E3RqWyif9on7OZIb5ERrs3YZNrH8P3332Kn
bEOn7p9nQ00uTVaKp+/Ui8uuJPmJD0NvAgqHJLjGZWTHFSKCHxO7h5U4Sg2LZ/YmyYGfbLRsqsu8
QS4W0mbHddjPCfnly2lPCVle8PT5l8cyMoQZ+X6GmxT4UjrW2mNqx9N1Cr8/3FBAEq0SYUT2tgS+
4M87tt/D0sjqfD3JTaPkw9pzcefusmvbcTvxTG6jM+1f5N5A0lMhjdE0lpq9ILGkPiwBily9BzlS
YExURtFdj3SiMM10sOISgRSDwGrMFAicJ5MzSkqf6sTxX8P2LJzEbBpSgBHgKWgxnZiLbCnMoaYJ
Z95WO0FG6GHBDF6/xOqbL8/CVNWiLeaNgwV1xCqqEptoqSO7UOkf7crVC8tUP91CFCGU6ncLwO4J
jOedWdbPXwYkIv9TORiihHVHsVeEyASLJwd6uFyn/J7InJHHp1j5dbbiRqQFv1FUNpVplnhI8uK6
8X4hCWPhcMxCZLd/RHiW8IHF2p19ey5vL4OZqz6CE95wPO99g50sBxTDGmiDmXNTsV3Y43A3VCDh
0BDKoeDV4Nt2bZQ4G/PfTU6eOd5655R6RIaHZy8ILmPp0zOxByw+jOTcEmu/+01pfE+fkDmt58MO
j74nIipOnLSExyvz+jdrvc4Mc2eHvPgd3jbGTwiZfSnpclDrimmzbtbyjW5Dn/sj02hq1V9Kt/7e
ThhdnoFURDn17xX+zBzNGD/6f4yFYSo5eyWiBSwvhY8Mr03EjGHqdI0ZZqYKU4VqpbrF92HN1hDh
fGG4mHV8Cdkvqt2sB6MV33J4by26cklxkpqOIBof29wGqP808tSUSxriqQqIOO/9VVQHuCWHhiG3
NZSpv63QuuHJUDHsNFqdxIMpOxbW1gI44nvis0igvR6d1O+VlW1EQbdJiQ2nZyKodmNV3Y3A4nVM
MUB5vRLO1fZ9rTWMcTRScMozwdy+EGrChWO/JliV1473gvLAeCz8YdanTOOxwaJNUZ/PdxREZNZZ
yl7OgjEKU3E/3Ieiha3pNrhZGeJDv8KGe9Z/d5ofnX/y7lIRQEbKTYpybHwAFo8/6RODbHpPJjCb
wMQ4kaZIRIIpDFcruBvL3rD9zCYI45jterA0I9hLS1p7q4kkKp5fLoZcpuoSsOgt/jLFQqekvHJn
CLgYWJSDYiqQJVv/1HmFKHnTAlsYPo0pORSELQasRD+FUFlp7wb0DR7MHxkmbv1v0UhRRuI5hXI9
rCUyEdvqHMQkf2DsTxa5SqFoY7W3f7OgYkqUGWAYwBVoVx0YlIoVrwq3UaFfpnAPNcPLzE5Nyc9s
nx2Lu1nAEBu92QExgPjI/+TnltJ1yoDZIeVjCSiH+LTA80ROzBzse8F5+uK9zuKFqNXrks2rvHjf
ZduZ16w2ukN2r6imudt7ZAn1luRrRFOr9dsCOvf67Eslc/LjgszGnl9bV1+s810GA7DAP6EekWDm
eWRDinNfvKRmPNB5rPm9hBJZL0AyiaFEMM+aCkWovs6DTIERtYK3yh+BU1Jp7XaDNrmABVzrvNtr
DP55hX8KeoNnMWhuzNwLA2+/bXbP1E2dHZMNz8BfY/R+MAd/lzM8pGghQZbjBwpIWCF9LgrvRWyh
clH3kNPK0xKsBuJpyZ6n2WHNS+rR7DbX/+B+kcZlb7Qj34i9ICQ0dQ8OfTFgIcXcoqM7tSsvFG30
gdlp8PtED0hm99STkjZ7HtCNuuBHuUuTm1t97ANxWptfSOk/VGAj6DtRmgFbJ9nXvKq8vOFiBr6e
8cVBnNwa9mAa0sSLH1uVjGXu3IBzykjrwYImfYFWl02RDc6IXSKpOFN0OH37n9LOOGYv4P5+EmZN
UvArNQezzuN2HFlngFtD+JwY2fS9xL+33plXs04NzR4ZaZLV7OHzmja13vISPVUdyF0Ie7+XJBpr
fCoEuOv35fduP6K92nhCVPpxrRaDfLOxjJBFQctvh7pt2vuWFqWn2PnKKn2Fapk3Qzez/JV8U3R4
AHTByI4Su8BDHI5gDYZptkLAFo6u2sPjKu58nSL+wYfP6rVVnLR4nNq5Als5d6CdW9ZtFj/CtYGf
w0cRmzwMS63zT2qnalxRLU7LXCLQdu4HvMkgJcXzDC1kFZaDBL3YRGm/dg0InyXhnAFPwRANjA86
glyWX5fvur1y6gVH3w6YjYtMRvuef1n50bmgxcrzzioyww7MYDO9APCU0q/BkbyxP56jRCd1AoFX
T9xAeP110SmbNSXFKMqvozf7bwRWNeu46v9ht85IdQrS4dLIW15bP0HRY27/fgVYGXK1Xzb8Mopw
4QOXOleGPxOQ4Drf38TvBlJEfVmGwF+bOlsM078pNfaAcJOqejv6NREFfwq/nkn00mWbqalVaw1X
FW+QmbVDogLJvHKfa6b4WlIMvi8moJF8ssZCne8G/94sGFiDf39w8Ayme6vqAjSUja99q0R4DJZt
SkxQiar8VmmJCXp5SXi9eN+Q/krvmCdA2uq63RRKbgTyShWeNv7o8OPFIZVnoFa8CJ1RTEfKejnG
SfkCuYeSRMEIPD2e7cX2eezSwcMpiSJDpahOM5EF1auCkQEm/aUbv8zrijC/dKut5P5mlgkhIHQ2
CuK9gUs9w36E9W1IahSuxKRfypLDErkaMnm7iU2jhvZnRkIX4df8c/Dg7HwG2M7Q7FY75TwIeQ4C
+ephjkQZih+1nc3pvO4c3TP+bEKy8dGuv75Z08T23d+lknKNrXEqSMGiNOI69EcO+DOwf0cA3Xqn
Mco5AVX+djo+qh5LIwofEBwl2lNhwPZk9sfSc9tvK/FPYTo80QrJf1C/SPf6/BgdurEy1hNONp/B
wU0EFOnOD5Znjhi8U9MVXhx+GV44kwQGViFerGsqeVRQm62NlRtNkcwd9pDWBJuwXSU7wh/KrFcI
qzW9GG8JGwtOP4bSFg8Kxw7NKGBs3sMtGf3VDqDA9/AQQbW7Qc0xnnws3lBlTYeEAVW5KJGWI3cP
k8kagKwcfVBeWCE4nQAlLd/MuwQ+kEZ+NSc3jqWrn9GUlhvBr898PYQRzN1Xzdn8hh79ildVk3SD
4NVi9fLVx92E2OaebXfRCQSNxJG41SCfHC0kw21vwxyHc39IKlDJBK+6n+fny7vvgu/N1MvsyLrv
dIDe+qfRq0eZAa6pzlbYDaHra+QEyFSnQqEkk3JztcNNVgTL6DJrnZTYF2GU1q3tXdrq6o8Areaj
SXp+6sRfjFuT3KU+zhnvUgqSt4e0xK2njbSf1vMbdDMBBAx3pT5limAOuyJU579AQael6UxJGTsm
jynPMr3BQXsm3y+zVuMgk2Pb7W56lnSJn8kXnoMYnT4hm6VUNHOMHK3bjjGLAbz2ceRc+DhGDF1j
GV5HQ/oc3kv3OsBJFto5m8fxmUxUmS8/ho0efWY5NzvUYr1W9KEuTok//ubQRYw1AF9+eM1Cl1Lb
foJyleEnY51Lj1JdIpwPYkEzsfNP2F/8BItPQm8wSpL0A5gN78EeVjOUzTeLxl4h1SEkyVpYdhyn
JtJczb1M29jUUeCNMD15w2XD//26iXa42GeRgq4GBWpMJBVhixEk9AJPKSiAN4n9K+UG0AXz9r+L
byAStKgud/jmYurcuM1GOrjMbmD5GHFFq31Duq3cPYs58Glf3/OWR2+NHQVKSxD+RpwAgGvTVRah
x7BzU5SfMPDg5qzuFTd6ypNjksE23QN5+ChGs3yxM8CMTMwMhNlFv8lnCxYqtrJSwJl6mR+I0Jvp
HBJvx877J0oUR9zF+xcybhjCNSBIRk4Nk8UQJ2ogMef4ZT70KIukcHwAAH4MRgyR2ADmiuxWCGGA
EKxtTiSyWj0KkskoS9H+0GXD9Bjuua0mJgUn6wot0neAzKWNxkDT7mbMuThcsipMganbruOh7XEe
s98lVmI/Kt0qNj3GDdrguQ/lGi/6eiSzbAqLDzKSuikyg1htboTcNarCHSeDAP2mDsd2dSXi0UhR
4Z24hr8wruo3vVhrh+5rr/eq1P4O7QvHTPuTwHLii4xkD8WSm32yI6YnHCXL/QEl+B8ou7DEFWzr
L70AgoTqpjpFyVCSXZGLS6T7UArst3JEqOsKu34HFMN+osW/U6tkuPzKpXT8yoScKJJ/PK0X9Yhe
xOoexMd8x5T+81S4CXunthvmbQovDV4epEZceFqANQw5x8uFRb/SnfM5gvOVTGvTlTj9VjLh/KHW
tefrTXMPSP46wfBx4qR1z93fhBLFWwAitqypwQS2It1c0nwISvEjo+Dd2oB13YyvMUUVRon+ICZw
63wDrTMpqjdaOcFfIfbUM6bZOR2LBW5DKmEhaiZ/dtY83e5BkWth8zhaYPklsbDPDMRDFalIhfmY
zEBfwp4rDsvgOUftGcE5axpaEU0XeE/IUwhSThwtW/QE0ZeGYl499wKl6JwgK2J3zedCOb7nBkpY
YXF+rgQeLP4ZvUZAr9WgUXf7mdl0o5In24H1OG4V9CjaxS0NAF1gRxTg7zE+6FTBjak1pz29aJh2
SMQliFPGG5fj9ucl1cInCSZVLzzqH4TVXD/rrLkR5Ax0mo4ubHFSLkAHxhzk5UXtDJAFbNilmmlD
nmQ/c6hV0aPfroh5TJxMpcBB3hAZSAULi9bT+nlVxCfiOS5k8OGvMSgiiMVfJvivLTvwaIq2ki5l
grQi/MTxTTN1VehkmIMigKphBVZWjrsN0Fg+tMn5f+wKJDDCy79bgki9B52CWfCd/UnX8Ps2XaVa
ofyYKqnxnVpSz/CbLbBw7ue1EPUWFnZEDi6kudx5FBgMGQrri4sj0duOtOcKk2FH4ef31iXqwsR9
9T+bE0in4vWuRJOpf9PDM1BAV9VhrknnyRF5vX5Uwac47UA1+MfWdA79l4mOIC2wJbmXbUWcpkUy
LRUunkSVXw+9O/kfTWJ6JckytGSkdzJjg0QK2zx5T0MlBFd61UfiwABUKNyq46CyW0n4a76bT4qk
Xg1NYQHqxa8Um+zwH9sfaqqsKhF1PRD9mEjRuhsFofdSRfOQ7pw9U1Nfk2KtTm0W5bl9MnkBt714
E+/jlxtx0h6SF8TM6r10uN+XFwmbZ3DQgz9Ubk9LtT/FXarDpJIocwZN379SvOaEEU2HJ0COjBBO
vwv+CC2/c+Ns63lrHtHbOd7TDz5lqT++x8eLGVMNdnnmtH5SuWFbYQFaUQd33jQVIc1SOITI+Kuj
EKCj2mTxiKcr8cySTtu/wPfvhEvlRBxy5wHtV59bAMkRzfRKXbOEcq4NwgSpZCNQY9cGeTkGA1c9
nAOykRv9nvGR8AlGrs5qS6LWybcXFD7rRJFWeSyUy6Z+ZHldA7qnRMLYnGZUtS02GDIAzTBXk0XU
F4yn7kH3bjhuOq+CnlCBfS8MNBrxjoocfh6lthqhhqaSQgFfuEyBTyJeaWXO4DdSkyuKa7fx3v4I
wJ/0IjLSggwH2T2EiEia5Tvus3dqiaJtBm1USG0XgMVEu2CEiJc8O/7Gjag6cx3Q1tRKfzAe/JxX
568FS5WHWfawVgIZ+jqwh1kzqbZMaShrgiJ36gKZyrd042mLvpNXydxnb2JI7krUq2Y1u1Vu0TRV
Adneh8MdI7iT6JRvfOgEAIw/M7AkFZqePCVo56mKe+a4K53zrC6n6QqVn+rE0fUbe0uStqUeQP6c
lNwGpagGFnVkqNz7SLA02dqpJENMxfcFU27LDB3wZ+2nRVObCWVMB+0T+yt99T0yTTtXlDLhEyOl
kpslL475W/mMl7HW3lZ4c8OtdI0qvC99ZIPSzf++SStJ3Ht1lfoXHffz2zqj/94vIAKmeUVETSAj
0iNkQEXJthCUazwooe56ma0E1645d3YAIs3GC3jT/gKK+f1r0qlAol2E+Z6+jl0Shl0c6JUUV0r2
cW9FDzxa88/5tqimaKTWX9ToV4vmTwsIUh7uopoGX4uEbqru55bvNrah9DLe5L2iGQwdEo0kZ19z
fqzx/pMGPb2/wbZE8+dKDnsG2qoRH8k0a4rmupSEeKmp0PrgdaAuIwZT0mDCBQSmviFLOgsr1HM4
pep/CVAIW8kGtC0e0t+DoRbIX08gL8LcFC+8JgyH+9IpSDajYYj06dz9h1XSM/3JEXolQTlPAj8v
y4n+imWmHzd7VFQcwTMcIiW6np53FqH9hqgMjlffOpH+nTyPfzFMg8itw1mqFh0qRyNDlyZHMNH8
/DBme8Ujq3suLbgutlCiRVP85WCF/NMPl1p4hpOzu9kY4J9nFhJEyjUm8OLcDWs+u7Ym/Nov8Bgy
JR/EZzBD9iWQCjl2gMbOwXbAoL8JRkC4YcWnC45nQ9Oh9RUWBc82oqsbUUsM5nJEH4NAket5r2bG
r2Ll+JTiV20okOQ8Y9F2V2agMbWxY5EIrNuopKK2mtVYE9sEGoNJo5/82YMCbi2yiwqwC21cDkV6
P26b4/YSzAUEmYGr0Z2k6VO9IeNT5EwZzBuNKINyD4uXhSEjNJuzuMZAwelY1dMrvchqHifbSY7R
uqBJ59714vaVeASb3SulQmdk4Eo1hfwvHsXcQClMIlkzqluv2sZSZq3I+cBGngFuwASrFAV1mVWo
qMburYM80IHp6rGzjVsCnycCBjs2AzHBkqQWUUVPV0zgZGNMcCELnQMzjRD2nFJOADiXimcZy+3R
dSf+sWSoF1LUdYAo4zX0KHAdtINW/4sPiJWLmmCnqemBuEERGnP9fCOknZ1/+CU43iwpEgivrmpp
B5PjGUVEBBvQ7Ir92QbYOk1u8b00auunjkSbYlTW5747Xza1tXtHjP+iGEuZNcr5RwaMvnmfMCtn
mZG7e9qeu2hOy+g4tuAewuxDhHQ3d1V6V3/DwmD8p9FoENWEC/OBt9L7S5LBX9nLhxNJizBdi69J
5UImCChfvCL4mdUxqEFcBFRI9A3euZx6ZVel52IZLnettP0BX/6BOMkj4wUc7lnPstDr/iW2KuQ7
JknX4zjZWxsp988EHhJ9xYSjgwXLcqiCOWiOU7m8pSFy2ZO7eB/dD9/1uVSE1Fr+bA54JJZhi00E
Qx2W5W697GuxUMWYS+DMYZNhBMLCrc9JoWr51LAK0xrntM5Ka0+kv/i0ysBcbApLglxRFvaULhXN
M4rU1jaADH5XMH2VU0OTDjAZgYhWkT0Obpba0XY3qS0FBs8GXCesUppABG234rNaWI+1FpaSIqzK
M5YzoMQ7vP9U1LWpoZU963tIS+vIGWIeudLtoD+ckvxsgx2gdHirQJKWeIiUldF0HCE0VKKqAFY9
tgoBtfG/JEapI+ThKc7NFzQR7kkITpTgeym5TFlIcmzDiYFhOiemJA37apAtqBVOaDMhugD4fVww
gGxzs8/FK4c+aiOSBVMs0iqwQageVcdzgoBFtcxSYntlikJdMv6m5jt7SP6M0e3ujJnMUhiI4Pie
QvCqO10B665K0oLqtn/jSw9z2WppjdDGXz6bv+fNhtRJuRml12Ui46c/C+2ilBKviFFzDAXgg7J2
7g1tfrdDHRPEAapnTXp/iRMi7fgYDsxbzb1j4i2rk8f5S/Jng5B+rL0gRXgPr+e9ymd2EWaiPNz5
+wSjXMO9UpLB2yhhua6LZdEZwIXKW+3T370Z5hwPUapbaODzpS+jt/S24zdTmwRIpOQIhgtD/63l
CW33iG8iUeELADEw4d7hugTWIznrjzvcd7OtO4LI696sIxYRqupTW5Iy8/NMbzRGbjgd8ZaSTcDM
ZfzMdR8E0RgJCiM5nQ30agddAIuqYod5/2KtMz1KuqksO31B3VBV3tH5kuF4sga2owkx1bkCr5vz
G4VOwqSHGNw+kTb9Nd+LmFHsnLBJ9tilpGeukScEw+aSVkzAWBHM8FvQwv6O5Og3VvC26wzvwHZl
wlDGZcgV7TyLD0mlAGNrGY6if4sjCrKNHuPdGnUhoHKA44DNk7R6AxDZ1VyphmGE+U0A9tZJ/N/W
wgm6iYfcUp7JknBmN2E+kU8kCzD2ztMCGAzaxZzRdKee3EvU9Pdk2ZYB0e+23mUEY3T/y8Pn3Fzr
FjC2ZxDDToTDHjU+Q6AuNHrFlVFx7IdyCDr1CLkmjDegfzMjsFKYpIHdUCMP26dpUa4fG/2aHObb
XtU+LBs4jOUJq96W0Upzegw/OcBvnHjT8MI13r6rD9JvcWK1qDuJLl/iYK7FTSEbfqTmT0FvM8zJ
58d6HFHYcfGkyYxEAjGw4dJg0SSFCX9gKyRb8D+N5q0zmP4cf90FhQdzncX5W0lgrVe3tOWWVguj
sEHryEwvYGheolHaJrMXceXyTXaf924174JwKzCyPFWnA68CIqLdIHTxMS2JBIwG0DhOLP1rNcvW
mOyYbZqUjKc8aOGOGdXFYkCfOgt1CZYc478/60ixwDjufjLIKEIONxG2cGqo+ODe6GiPmqH0cApJ
r+QJ6u8yd1GGcUggm81sOMacneoRXtpNYrYcoF/YkWDnfodfDe47oFt41BIganPSF0HWLNTXuZ6p
gaKHZPhPOai6BeHipbyZFpCFzxAlbvQEePW7O95/14xiqJ+rXKoGKE3+2YRRYYCMGiuEyhwc0fuJ
ri7pgx6d1x2yPo20fALcCRZ2wv7zpnaryq/qSrXuQE1+UfcUmxZrSQoTPRGrk1JMp6Z7IkYx0qMf
wFSep/XmRMxBtBJhJD6j8x8gtuclPi2ejoeRDhly3lpHbMYkPsNrF//DuxRJQl6hggElU13FHg2D
ymW+zdcKmtziuQwh41DeUayYhP1C/FrH8XTupiSOj2ZXj3ALR7tnH3NmHe347vNEdFMqjswa8W80
OUf6kzcC3Bt+jNnudE4cNL23NujIGFms4pu/UWtR1DSsNymEQhqcpiQnzjzFgHsG3WTcvX4ful/u
BKRSMfWkajJD15tnI5IgBdelO948ruudtlJuLOdq23ZMwpdu/b0XJuJnbypYh+iPCs8mZdxpv085
I6BoC6hVFD8QDGYyWWEIHRYNKy+10g0wlrKIXmWANLtlsItuUCaQqvTdC6yPYcPwtmctrZBXf+mf
LK5Wf1Zse73i09+0uUyWKJ9QHEoervb7ftfeYLf6RYcI+v3zJN8wZBus6xHit/cYoQhyO7yopqvd
3Y4stsQLR1YywywQ2XCdXWbWy0CpOmshfXGzm93/4giEL7VmegMrGUeDLkguZxJ3Ok8jUgVJCtlD
a0PF/VWWh6E2olXbqPoeCOMSr2O8ijsciDhXCNFCQyys4RWyxw887idZ3PuL3ewJFZhBrZ1z5dVH
MpVwf/BWkBAbOZFhcT/Is53+YZEII9o/AV6Yny7sk9LpIIU5YCmDFqXQYUuuFiWMvZeNepdRbKKo
ELXmTzajflKD6CvaFKQ+j9JFASbPs5vkMI77Smq33rrFR0uUfHj+PTsumM8OG+rBcDjwowRhEtzJ
l69wnKzZEH5HwE0pOGjLdR7oUN9rtIdcltUBcaJy9Wz/lGQ/+svfMBEg1dZUx/Cw76zRU9Kzm7j3
YFClPS1GH3lUDRwn4DnsXuEI64lTOdxy5P4kiL7HJDkeEkdUv77bVTXR9ApLEQO/pkYWGpQEzHV/
XTdyM1cJbAVbCLFVTouVjXzPRXcfhhPDvv15UQPMkmDWHaZij/K2NPSVv8Z3Ty8njW7w8m61FHK9
mZUkedY8lV2TAI4M3vPH2mzlv422N3bCKDT4KfJ7iUfo/NMcauQwELnN2M8acXwIxdzN7SXKv+sU
AQrHxVAqQtkhAOHc74cXM8IC/BQmE0fcbcvmrcXWQpP/nLqV2hOa0laog6aUZRIjywCUwPy5MWVx
3ItbUACqQQ6bCoZWibk4DKTo/Ai33/GrVbwbhNWlPSSI7zN5jS/n/ZwvkPaY1rCuuugpA9Pgia+N
XWBlpnkgqLBGXo/xLrbJtVpX0M9dPtHos+wzoUnDFFfMmzJk6SbW1EtOORir1WMBEuH0x0tUVODM
ufqFPz7aVrpujoCeOTafBceuesFASVJdkaSRG2m1V1XM1CYgfnF2vaw9C74j8Du3sicRZTw/yvkn
oXEwH9PjC7mB+Va+h2f/jqXmqOWjsWYyKzmcejiYDcwiXWH5ujBJSLMLXre0mLRNDEc0S+kkYJmI
2baNhg76p9OGwTDw3/7YBQsGpGEx1+0Wcmkv0cKM8apfRlaHfE1CrYi9w7iOSZoh52CVDTBVGOAD
HzM9SCN7kzXKGJrim+Ls6Ml1SA1p4uucHGQ1QwKzqxuzXQUCkq0Pa1G1471y84Os8+8d1lzgry9H
e2as0Hh1XqA+EWOHo04KSlNAyvdze0mD7PC44ZJ97pKRyMPs4s4PhRqVfDWlFbrxCNNdbUI0dpF2
Tq5BHWTgfvqrD7fsbjQFBrz3Vdnw0J/ERoiIOMK3JyxfPbDy1Zz0GmBjL/VIsUpqmKpxtL+hJjsh
lmPjgO8q1vbopZqqdU8WZKH4kq1jRDy4opQNv7N/tVFk13qQHt68ssNlhiBpqlhkltyUA7mm7EIZ
mSFe0GiSok2i0bEzBqFw5XkXdTFvlTBkOLeCvshgRxb4hDAtG0zzYU+Z+qLCcnPOzKzZm0hYmaEr
s/wYcH60U53FcI/oMqxXpyGpAgPQh58WM3Nn7tLJ9HMyK6yiCxUUGr4CIYPeUJLXJd9zS7T9zCaS
phvqZl4CuubpePdw4dclHvlKa7h8Pcc/oZIO8MH023YjxzCz8KWzrpQyGSca1W6JS1zZvng2FeBS
Gi4nE/1Cj78nRuMDOJmTlhbhoovRBOo5YGF4m6UYcZR0RosR/4BjFgE3ek7w/4gGcr0xTGNTdK+1
sJw4UEaH6xV834etnAD2/9XNRj0M+uZtvG1NtxWYak+QxrsN/KuzlEINsvo83Gm6ktSUXhXQ5bMF
614DeD/M7ZIzMWNsIJjsEQdh2zHT1MTIniP8SFB2FjwFG7pWB/lshPAKMXJrCUIqx2FpVee3C05M
Zt1V9reZCSCZCxLBkBIOw9ZNtb5d5syjYSfwABjGQRVbiq7R5ItgRo2hnWhTSuCI0babY1ag3Vnv
TRfM7Rb/y3jdtP4D4E+Sf/g+H+FADElnYZ08b6sVA5swCNSCqvKeAExDx1KoOp5yICD17i4Lbhnn
k8P6r9VxCEpBBPBgCazenJ7pW89x4qeRYR2Z1u8X1Ose5PPwudHOXoekJVt4MIl3VPHxP/HoDytL
5i5QiAZNrN9ffLBGrTcg9hjgDncS4fBR0zIx0aXD+xYimoWze0jWyiqWP8E9mEdMttnjdB8TvnaW
Rnxcrx/YxvQ3e5oeFsxOoM2NXDGynu92yqbUzto0kjq79UmrPZvU6m/v/mS1Fbt+pK8QuVjTJZbH
5XzhGE20mMggzEFEFeYPGwqgVh8ain9BpnFCE7eUyB0UxQcQ8S9YqpQfMTUA14ivqCzjjBe5eh+J
7OTR8oKheDJnIqukrNnrrrrCfRFRNVZBnilB5h4ZIbwyyAAVlb8zQQND5ZnQDVnpbIsusZgc5ElG
jornUtD6kbr+Bh4vt+WepTvTarxct+QM2nJZdZSEiYN89tz0kmVVUAOBrp27FMHttegQ7Q4vLt8g
WlzFglWACpE8mylQrVoL+/soWDA/xjF/GMRlI+Tb4uu8qbhuet6mpxwYwQJMCEjeW6+mp2aUyL6s
OE2/Trc1aYeO7xm+Jy0uQcQX40w7fooV4CKMMowiBNfzzbfRrMALGdChw5ltnBkshhFlbx9IhB+B
n5sW0EK7jblUtnIY0gKcbTLiwOH7yboXkiwvVnpq1LQsp9A7FjPfBp1mjAduNzi76cAYZCmnKxCi
2VNhIvPlD2NyIYUIm6r7YINL06H3IUVkaVxeSHlj2oT/U6Bw64HsTBQ0aB8pQOXBuO2Tv2VGWAjc
Kam9mFy7NiMASV7zOmyH4Xh1N4dBOFGybzJxHmkJC2bZuy1/np7ZEBJMIyusQTM5DSTZQ5WPHHSt
WDu5s/bzVREVpvEmcP3piSdAMynOZ0BbJ0bykWy5YrIGe9reNHQdBJmNv1w6ctlrMX13NpaJBDoY
YjepeHsL1Ucj8H1vCcBRT9/Eh/o8kx5sYP6ixoSlS70jb526eAu4KHPvKS9JC9OqHcFjf/ATivHF
jfDxCRfXIoIx3l9bE65l7OXqCF2M2/xvr1l3k9WM/YsS9O+1ni0gUxueX/SSSP/eYt79c70kFo0Q
oKMg4lp/nY16QKM8aBrn8r8t+zMErzsVmGC/hKHDU/RXBQ2o1FrH6+2rEMIzXz6liy6UyX1AO6R+
6hjO195d6n+yaMVxoCNjkqjfHwJoCc6gZpdrIDUEG60j12tWwA2oSs+Bluz0cPbQIdKqYFr3B2o4
FpkAcz0igXmwUU6v9CKb3mBRXuIdQZmju2kmeg1931d8Br5yv+nqsLdZaVFsy8zUYAePx6F5ZH/p
WZGA5uJK4uLdcXLTOrLkNjun7Tsk0wRUN4/3UJMbZoAbFbxJPGoWpIVbwz7BEXjXQYzucu3GWUJb
OuijQoHZdT+0+Q/RpbrWvnKSlBRnM+JQadc2fc0DDYHF2ZpYVSbUTQ8KKBn6mja93PPmxHpqLZjG
1ccm0uTMI2Oyf21qnouPOtrHm/AtnUaAt+vxC8K5FuN3OUVQ+74Q20RI5FLI03+lJYWPWbWjK3AU
FqY+uNpEv4ZlZL3aSz98AnR+ehgSzD6jY0Vje3i0K/WHGW2Jkqf/9PGZVjJir01jV3EvZuTBhBUY
NQoItvxrayKU908K9ERO7xxCYDH9gXPEypmTctLgVhTUe0h/ywBx7sSbr3jCGoC3oZn6rcW00pkO
/R6MHhevjrsb5bLu087xcMKJ7p+HrFlZ/gsZpI7VDGcIBjzPso+dHLy8iwaiEVHVWlKmQRnXkOXx
o6sxdzQViRjbJ4v+aLZEs+OUlvLIYig2WJX6kV7RR4DXJAMNosngcUbuAHDFqCOGvhibE/LLvpLu
lXHzsTJP/T1jawNEeXZC+1j4OiBoeK3dKDnB2yvcRaxNJlYod0nsuiMjlNa9yPgsbflE32PYNAce
vFuUQhuVVIr40UuPINp7oKzgV0CoSvWTfVnKR0gJVU+O19GVGQzQN5zhiVEypOGwou93qn0Clo6r
37WAIbNQPzYnTuT8oNSFaeXBBGDFdT/PvQqduT56kHhyAnwB5QNvFK/jX5YibkzG2SZ7HIkstQ2o
sCLH48Kh4gQkoyJrEjV+JU1uN70wJbL3FrOBok1kmYEXEx1YcZbcb75YqoyE04jJxhnolaCcpmFi
l2LzYVQ1XDPvGsZtQ+sla73610qnQztqbGORIthYoxB6HFJ0xQahJfOkeD+MQN8Er+NWYwmAihfm
BLXlpq8qkLK8pWu8dO+iEqL0BZiOpDp7IIjRQz9TaKuF1GIW32YZa+vbVCvwlfOwT3Iql1XNvZ5Z
vLSwmK6e4wbUuTU4iOq1tjljNZiRf1RZdjmrq2m31BviOhA+G2ieDqCah17wwNbDVh3USsk7PU1E
gjMCj7HqkN5Sstkd8S5vyuknTim0zgL5LJYhjzXBNlU3CusEx9Xj0Bq0Gx3wdyuZN5MYsbtEXIqn
svQqbehUAMYCzGHorY4AGyfWf1der5zY0e5K/ceSYWss9f6qFZtwUeY8Lw3y//rNQ3VjxzJ92/pi
J2D4A8t0epAsmKxR+vq+kjbpFakgbequEWH+iUiT5bD1ke0jrriR0WyYUXjlVrlpOl/cWCJljTOx
/5/BRm468+8C/wdZaMxuymm2H5rCCLw80qlAMKgy1lQaOIV8KdQLud+YjEIf3oOCVilk3oHTJJxo
IJwF0qMY/L68vRlF+/ZGLQYtfdRKaNbkg7XeQZP05tiHelTofXVl33XILPqUKkwyrQ12/wYilvh4
edMKUjx1HQpwVCCdnHv0qwPjMeWpLe4lRy3+21geSE6mKAxBtJ4oFdFvg/LuFgSshIizcXjmQ8qj
PmZRfEQjDL937rvwRuCBoN+vwodF9cXKCdZAlXJJB9OPRncPpr5PhANmYLaIJbKkarWCiqUyov86
fk5+EbrtAimLQObgV+48Zpj/3z0hq+eWFD9wdwtxh/zU53ip5Af3R7FuG3OioQYnTtZsFXb3R0Ns
6qRmfqM6LVCgBCO2tZrk3MYIOipPWzWoQk4Q1s/e5NsdG/eb6JJ1TXVr1ZV05QFo1PcEyASSY36x
lX4QXmQRtTB0k0vAIkSiffANSTyG2m98SFTlPyvbPrnkpPOCg/rexo4/p0fkVc+83dVelPubZ7PF
8KLnc6fx7iK0WXGrdRhJ3aMdRFX2Mo+dQ8+3SxqUsqGPZH8091oHTU4nYLQVt0RaEpJqYcxu3nWm
u+/Bd/cLLoT7S7DSMnhYcym42RJJBBSBRpK2bj5e9bXcAjwYAAf8QN99Gp8AxGYgMlHsxiLWAEC8
/LOb9ovSe3RDQQ1+za4znPzhjRPVkFqJ2bVIbFASmCNldy05olOaX39GrlVeChZbqujmN3pkr4q9
sR93f9LhNOWVmIW/Ybw674ciS3uIHrvJ9/rzyHWuLNJH03uKjZ0sqzMkrXmd/1BPEadSsiY4xpD0
j92IqF0iV0Nbxqs77FvTqBvfB/aMoquywfrS0y9AbZyhAztNiMyFyN6HYtwHkSq0s/C3kQd6qMDO
8VujcYx17aaJapbCYv8rrUIljeEO32nCWulgV/I3boDcdmZ0Fpw0arD+1/qzGvgTJ+nzSII1LXOa
y78k7cO0dS4hbZW/VsZf9mhvzBeU2kXzLjfszTTulZEIrZoTFY8x7cJH20xntQ76BehlM52ixwTi
aA8T0IZ7XizavtATCilpyrO1hRGBj4m9cNV5EJTvdu96NuLtzBqQ+5FJ4NGC5q7rDc3zHZjVIKys
TEynEYIQuvaPaLFPLkLrg1Entw3Yu5pEKoP41dJcN/KRRk32Nbb5CoUqSjPrxqW7M//lNK3BAP6g
oXggqWF/kEpMSyNSS4CsfrSTgF5GkY9Noag/dhNEWlYUUlcc5EQP8SraqrhJuX4jLvuQT9JwwVaF
70hL8UC8aGaGWxIkFNb7rjBNPfcHkJeLd6TjOyUstlYnGdyfXrvBVuEAvbdrxlocCobR4o8XX2V3
MLtaDHXYuQmtHeFJm9v8wQJe+Qq3Viw4/oUnYEHbsPE56t4wVWFLBy5yQzbXoLIYx1QSCPGbjSSz
vUIOvKjwC9mlyjMq6Cs5T6/kJUpkV+zvMThtBsuhQI36oRwGv9tchynVgVRt0v6P6boWxvRd/PTP
AkDehGpYRcY2/DnYS785rP1Vd6bheXM3nd4j01V9153TrAZFY5DJ1YatTLQ0aM4hhjm4tekrD1pM
kJu3IEegbVXUX4DcL7dN2WkdYOugRWqPJuh8TxKz1V4Ef8xdEByDoZWVc4sc/mBtYy+gw2LW8VNL
X0UoqrJz+xEJv1kxhzW8ErvYZQ2nBhkEzHm+DionVHHNJke76r6cgv7X0tjY+fk68+JeLF4SjF1W
2Zjz6B7Zfv+O2dLcUQj0DBz4JVEU6KSs7Yne9EMNw4nPGIIi4PZq152N+vdl8uv54D2MYPmsXH71
C7mETpY78CEl7FavEsEDbqPqCcFVFebqj06NfYE2P5ZWN2ueUbLaDEJHS+S/cgNA+hpLUtNaqxDA
IrDC4QoSHTHxgDcelfsybFJUIJSfeec/xNBVfKRF3IQU3YWtIfiq9Nxm3VmP1ALn3CYI/Z326Ny+
MVNDcQZGUKB3gCkFMktaVcSVQF8zp4S8ka2mBO4VKFn1Vv7XY1LFQqdWqyGrmK8nuSYZdqRGWhih
BUwQg8pY5oowbidsiclDBqzwDHK7wuSNrkk3eBbQLAMOSEE3sEHWkhB87IhcDFT1O0Uh+FRJVKqH
IIedg935+z4Z3wixQJt/nm7FKTKdyXl/fMkHpLB9dpWNTtiFM6gjU2/41DRbeh8Sj8rxLeamQ3SO
CkeEv0YgSfo2P9rwhyfDnLQzsPQf4rBwgJb3ROOcsFExuPHMeUfiGhkHfNJIJtMe3TVn5dG+9zIb
z0k+JH3nE5NcknvqZIPEjK4S1iS5XAs3cmrrbdhZ7ziTPc+rgKza2dxcjUptF+aNMu6l2Z7Wp2VZ
tu+fYXTs7C3ZotbvaqFDei2B4ZQP9Sa1OAd/9c014t+4893zRNBphFYSxkJsJu0/m7lrqWeoMv7J
gYs6hDQxad0c0ZM0PvFXlko1lXoOubaIPMTN7cFng3U2ky/A4fXY9ZR6OoPVXpofknYoVvr2BAr2
3QYXlgUI9Z4/2LTJtUrlM473RN4I5BIib+FjtWFWgWXvFRTiogBO5At2+wEGpX3LSqQ+g6pAaJHu
HShcPRbiY6ROB7tdgeCfEsT09c5Jnhcp6esyzPA7tRcZn7NkGX2RoPFEo7S6oa5J6MR/SCnJuzuT
UFkKcpnS2U+J8pUfc4DZ8v5fuMBwnh0LA8skxG+PQ6YwNh+2I8W3r/FaEIApkFJSvm8s4EEnTwME
YPOFwMIkPTcUo44gcmYi7UxNPJQTa7uM5mnj3Qg/bwR3PKMhKGKnZed1iuwoYayyhO5g1PuhzJNM
RrErkermXEzFt6S+NPpqupjK13zhlfvsC+MM6ngULLgAQpskO9Is5qf0lcIn8f3fmAPzq1Q0nBNt
EJMIFm+O7EfOyAaaxdC1vF/LIbkExa8ZCS0ubvNDhaqVMKcAf/OnpvSBdDO6WM+lmXkIq1eoHBIa
0iiL92GHcF8xcXjBFBBbYjq76ZxGsKRhKqyAWUz7DKVAOGOzLmLPc5fHbq9Bk9Zdo8Dc6XPbmxCa
kYxfRmOsVJ0IPJUZKOzQ8O5wDsHFyZhYBswKwU3vUH0G0Im55xWeVVZRhDjl+rdBKCB87JOUB9Cg
a4JezPBdWxWNrs3cney3xfbOEFFVZH+8XSaPouT151miJtG32NwIgvvVNgdMkIMNEmmg81aaVYMk
b77H9l2PkOGwD46xqaOYTlW8vf4goYTpK+5QlGpQAArZTspaGC6g/a7orJbhsVWGM/vunZBxPUr9
OXggdyR6De11za6uvEeHHE8o0oO4R0pkquQiKim/7OcfovBvAqTf555vga6ewec+2iilGLBHBGVc
Fv/nofku6I/+dAaXf47zu+gaJ6JJ7lSq13UaYWP1Njj71CvfKg2TOrPZmGAq6S5BrIhDkmZZnYmO
cFg62BvfcKuD4Vh44J8F9vtOGOTOLBCReaX6T5qoujoq1Z8w7Pc8ZUcHr3iByHP/8TitD+p1mlb+
GC0X+CINXkcTtOndiMIYMTD9PAOa4Qygo3oZmSKdqDID5h5Y72Iv17CR5vTl8TFpaAMOymoR2/S8
hTmKxtpR9lyCtUw7rq2ibCn1F3twtoUwkBBpBIJ6GlYjAK4KLmZp76YU/dbotEQLdvPY8+18zCL8
ehPnSvUKpp+jLjpinExCBmIeE4ogCtINNMyA03niwOCZ1p0Dd7t+WqpKYFGqMV2+O5yDd1sbueEb
QedolnXHgRiGjT/McwoTyRcQZHS8t6WPpvquR1vdymuCpgjQfxjQ9d/wMgdi7PsxwZpDh02xCj6P
zu0dD82gS8Rmy+hqEvow6FpBlrNSvcR4hc0JlTaWX3b9Ty+wTmZe42UnxUjqORx7iCfJbGiXwbR6
3naodAi4HI7+594ZymkOKkmpBbsc+voyDzQenMMKdPoesNrkeZ69KsoMftkSRtjC1yF6xx8+ct/O
y7FtjywtesQ5vJI4fmYtOHZwOyH+6XOo0q1v0QV3G619Ejo92AuwE/D+BgzXkbtoCT6zBGA+uIdZ
N0gABUH1fRIVDnlsC3ZfuxtzVtT6dtEbMu9nMPsgQz41e7Kl5nkdEdHqisPwLXp1zi2cxkgPnbNR
lxOqGPT9qiYiUmRCFO6gqQsCSF0ynbQLTNaP0A5JfjjpWTrH6vu74CFGg/b0U0ir9sTXZh5OJAHL
KbtjcDqNzEYCkxB96TVJDLXSaPDfAVZhvBbT3TO/HQbzhZ44nSZ2zHYKgLH+m3OeFkPLua27+smA
Mn7y0v8fl/QEmnB7xuP74osRl5wFPCB5YHJlyAG6cpZ3hhzxw4B9+9UvymSUktD5nxW1RZiAxgpX
shBFE6wHLBmaTwVjSUtDkX9TRuv/X05EdLkCescbavDvxxa5a8UCkb7W2zlcCqmGlndyXQ4N8krz
W1tZ5jOUoWHb63XtSpkNUEHpgDAPCWWCqtW3XyWfLGWu5T6ZHBDo4DZktUSWwpmYYp+9aVnQDepS
CN6jpm5oi7QuNLE0YfNbHb/cR2ETO3EvzKy2ukPbQbT1QfhBEqCTH47yOm1lbmiGp4f6lk/PG3J/
pL7IjgG9PSWU43TxG+4f6h0MUoKSsx0klbOswiVZw8WjUOpUk1bWh0Cfh4pa028qzhv/r/UluvMx
6xx/M/KUlIyQAuoEhNjxRpic2Ygv+qKK9ouUsyD3WLlMHU5Cweq/Zb4XOzLq1u6dNwls/3rTQ5vB
Hx9SlpQXvzlrUHJgPwONZLYEw1NKdR+cXLBTxd5y2jNV6VjQoMZl15egPDYQ1CmZF/Qk17TLYQ4c
Dq/pcM2QfaS6blNcDHhjzbBmbBk40sMTlhBOVkAv5AK0BsjbM397MPRZ3ACXl1WA/YOwIsYXYVaS
TYQd3XINHesyY7tb2njiHgEAh034gISbtiM3pduSlubTkPVGxwsskbgK55LDnjJKYxFYb4wgb9Lx
az9UX4S7TjZTq0AkUQ67U1SsLGj9X9+j36ltfLusGtET8Zj38tRboUGgHa9oUFDOoxkPY+TOl0fz
fnI4f8YUOkFXs1BnFJC3vdntxzT2wcXHqg0ZYazXT3ZqEg8gleh1lyMxZ8kmvgzG0fhBGUSwz27j
jQzAWkeUl7VhW/ixH8sAwMD6vPRd0r2ulAfns7hEbvfkKYOlej79e887wK6+ppe5gwhCT2ohjhC/
M4PDpjLPRW1W5wFF0V0O2iyzrmPNLJ8fbDYVWumXpF88zfFXNymUbeuRHc35L3/7PfdBe7Gu+TNT
wy5Ohe06dDNRQb3H+y0tuD+qzP/KGU8v6DO7HcWtObsYNj5saANlIUq4yAdyOqPwOHPVTnEaLJUH
oEKha5f2gQyvSjlhjovgn46Q6PX/Zjo2UNVmor95jwqJvfc7hMRjr75yBeICvGV1RKThm7EbJkm4
9XzRn2iu8Eut57wtc6lKqwAvCcsntM9CVUMihNE/QMvZQFamq/9IbQab9aazGpuWxs1zus/sBRF9
grcLS1jb6cDXfzofmkUkWPp5RC9Su3Rg48T681m/oSjsdpD/3VDKDEB3HFNPh+0UdTso8LZOJKOe
zT6n6PiqToZYh+HORo7Zp6L+Mn/Dk1QHPFXOmYvKM+qNskkEzYItzXIkDysuv5XfkeOZJJkp0vgK
wcNaYrCtnmZM/nzeVN0kWqCqqFLdF+VVwPVruvtMQJ1bPet6+Cp4uDlgPRA5VswQo+nDTyCgtu+f
nUDopWCS75tA+s0sMA++xahGn6w0N9fgYW/8xpGGu4zh8dNKPEoHE8/M5wBJyIZe7f4aRAxPA64+
bpqUFHmEWIggMDt3Cqgsn75iMyo+9VpNLe8PId64q+wbGGLDplfQbKLzMrU5z/gfjW6fyV/zFuod
9hRvwlxojgW7tj4/ZkOTx86+SK/bLA53HmjyFB7yxGMyUK9GfVxyEZCv5XF4iRmKiZXooyiZU6h+
W+EAj7IRt/PbfUnqZ5IqqGsXbC/vNQ6R2/guOmAfbTqiB3y5wuH++eikKIBo81qFP1x2Y0ycCyjR
C95Nj7sPwTW2Ewr3RjPSduIYaVBiNySJPc9GtQSbQj+cDVIZYtXuWoXSq5Ek3zLK/v/KzUr02j8C
gCy1ZCGTvGnrMqE0yGuF6O2iFx8KJo8AFqAqECgrxLbxdebjEBYYERoE9xduQX7SwE04aQD8S/m0
jh6v9A/8+1Nsq1fpCfSk4IrYxwpS71C4S9HhyhhX6MlVocsvOq8f0fB7Z4Dy4gyXIm3lh0GpRbnT
ZN2GcdLMoi/5I3dhM7s3RwwDcuvMTopMZFyZM48cEEBJANPlHi9VxADy916yA/0vQV7VwjrQA6TE
F6Z9Kl12jQvKnfo8wSTZT4AGKIzRiP9zUMjQIoGjKiDfgUPRXSpi5e2WkmpI+s8PsC3RNL38fhrv
kpbdK+gh87yHmnWebc7nBm7TugfKEefdn6nz3qw86Wz3k0bsabQMSA8ypIFNvY5nr59ucdB5Is7B
IMyVFkme0GRoykQvQLsM8/RwgZMgD4cPKpgNzbisyzA4HQz6jvjhHqa8do7qqiQGs6P7fJUE039k
o5dzMigHvpAWLvxZlG5To+BUk0qejNzjrAZs0fHvH+a1+dd7/Z9PaHj7HwgBrXHNU1o7YVx+o8bL
hSRH3d4nqOOVaC6XQFjkYtm36erXcJ5c93yoDmizHMP5FEpu+ayZBrvuUSzSxMa6ibkYf573mm/N
vcVUNOSfyMwzWHESUKrE/kz81oLA6nnQzecoQr9Y2AJtyL1EwfCjaOaS6xxsNW1bhCRgjd2u4aYM
ZQxuo15ka8QUMBs/C45RJ+gUQpvl8392Wkjgdo+WD1pxdEKassjUAeDUFTyvaN8S+EEPhSV1bhwT
dBLbg4s35wL/Qj5VfzEAKLeheUSOn+rCcdnHbg+CFgAO7mBaUV3aAqVOwHrqMGRvVL+FhU+NdNiP
/ZGF7CnfkisKBMxLFxXS21h9OQnJq67M+jBvaNPlUy8xE9qmOJaReKQ3G/QHq1KQPaKqwVi1r+5P
ItfQ+fejf/BP1TmT9NyL6WHsVx8yAa4Ovlpbwafl4XkNvpuIDnUOWQXMJrlRz+qJtLsYv0h3/Px9
TMurNTwm9p/IMEACT7SgH2uWnodXVyhUltLQJfPb7Ks/VgEqQSKXA3QaVnUukR9n74NGvJLIjU/U
035RGcnlqzGuWKtafJbgPkF8JHrdFgCpL2ScTKSutgx1trx2Y8e0s08/YrpAdLMzzraaiIDBcuaY
dAFhumjrdGr+zRh55TubE6B2kB2Px7Ypn5uvHJD5obDUlEDz2kX+2lTmf31itnHyCLKadVrx89xS
0YR2Yc9zTylHp+qM4Q4gYKp/TmJiogsgFI4HifTObSHMGWnyYEz6eNiXwWJ4bs8yHURwbHs9l7g4
dEXPDs4KOOOzjwGBKKpLAgoVp0hCrdeaEnOA8gIM/EFfoV3rbYQJyKB0kYQK1wDMS17pQSxdPkjY
wDPclDsjm8IJhPhXuzh0yH63+Df8HaoB+JxqCtdfs15vxJJuizNl5whFigxBWDkwKlyU06Q2Exj0
rDsfC2caK4BbG6/bAbpA3t+HjXblcJvRu76wz0/RH5ovnubABEX2cyO9PvdC7afJ9GVOtiItitvT
MeeQWO2Rf438ABhA606QzXpE+WngyExMVy3ixS9nrjvDw0ykz90dmr47r4cNYxD1QuN9eFdW9097
aDn3jB1hmOM1UNcAkJCJ+2/C78ltqCtRKGmxborPz5eRtuX14CcURBZiGV+/uupi9C7CwsXR/SIB
9nULC/NSyYhcpqzhUnsynJHYn8dB4/qsPkY0WSuc985NnaJG6tvNKe9M87SiOKY/vY9lb1tPaig6
layDvPKM5iO7+RZn3ssC2Pxtl8k/JDkINY656NfblbOytG+2KtDzPRHITWx0L8AB0UcMJGV+WZvv
Yq8RKI7Xw9TWbIyoW3OKtvUF2Kd4Kg1/ZdOz/epb2ZFJ9wtFOkaoK7Y5w/CrCNhIS9AhbG2gK/NX
Ve7pBU3y5fx6czbbbdZNhZ17xoaRVb5AK8+pCunO3Q9DXpu5p60lJlDlndjQ+hXq3D2ESkhB5vwr
NOQC2KigHox/eSyXoGqphdOoavN2lueQx0Rb72UtkYrZsw49QIkU/IvOD6gQsR840tSaBi+NyUh0
VNUpDNbPu/tqBWnD3oDKUXgKwOba/SK8BcYtPlk+JXWgYncgYgcQXGl5cGHkUpSw3ALGtgGgDqzC
XrtE+52kjLETG6KfwGVf5PSnumXABYTV5ZW0Gz6OEc4d34NDHVP82rNmUU0M7iNb/rT6w/Zg6m12
/Er+A3dWXJigiIUnFrSW1QMsoqvsuZC3zxfXqyn0lL1RAczymzkS4ffjwOQhKfDEKTM1iforA+d2
VyoLkWbK8FxMb5Ps2gR7v2NdV8B4Gi7n9bgzKLZChehx/IpYAxe0Rc1ATYRSx6jK0C2syw0pnOQ8
pgSzJxYXx5IZ/uxyZU65UC2mn1MESt0rr6RF1tXynoO762guaDxFQFfUwRgy9jOzKMx13p1oyTLP
FQO5L5/GdRvRPYW3snttVbBRYwSG+HB+Mp7P36M1FpCohDjZuvFsC/D3ueMMAOpr/Jd91g2kitME
QcXHUCuKv/XClAWtP5eG0f/p//9K+ZcAw/JQoooDh5k+d2GMFhuSh9ekeYqZj5EID0+u1ks9Bcgz
H4qMATH47aNVpnhnNvhrM3MDP2A/NstJYbDvcL2hIg6FuBuxJDDVKWFAuCcx12cJbx8m3eHc+BgM
jJC35Q27BhDYhHuO6zVRHtnI2EvX5MfQHJSvYnsp2yIVlRoHtVOBnRV6W6HI0/Acyf09es1YNdvy
u/0gAmNB+TqAraChXXeqAyKTdARKjMupC3Rx7FiN1x3rKxVGmma7n68i0OUulO3xmAnJRQ636szh
DuaNbqmxTDwaTHvR/sGEUrlL4QH/9Du2lEUI9LkWm9dHmsUZCkTGJ7m+EU69IEUsK4Dqxg9/P9z8
+e8pNI/kB6J8VFX85hz/FnYAhfNI0RrTHrzLEL97Whzjr6Ute7nTtt3OH44uzQRbk6oCl0Zrx3AQ
Z2kZjYQHVYY6BOf9u0/yLAXjSWmh2msp1J67yZnBCtGusLVr7SMnJ4MAdGz29AbqdNehS2ADK5cU
QhGmAa9RmPq2hnhD3wIEh2AZO8zV8wZ7UHl5b+PM5xd14FrpgrYA5WisOX0tCl40x5C4BkTwvuQ4
4/ww+zRQvBC1Cj4Hru+Vd0I3+voaCMfL/JlVdE7pQ6U2jWHQwBBluJJ1p/5vMZeRoPbmq/KTAksh
2n8sp/nJCfi0eLXWoo2jwngPexTPDt+gAH9nGhhjPt89aE44ZK7QplwmpgZVqpl1Zltn9gch5Wvs
MQ7zlNbgBsi8m3gaZPyUBNfE0SkCo6Ef4cC0Ftdr9w/n47fUkUdv848gj84Bwo+vuDdRSaQ+56ol
lFFSi+5iZ8TMXKg4Z7mnr85FGygbwiCWdGYPUK2zr9+7ZD6yKP3QC7S+jfeKHskEkl0v57yYltDF
kjRe4i0RFi2pIq2cAUIa3ekvJVTdM6NkmcuQBUoxX4+wj/0IVgdiRSWW07pj+jRRnX0SFztEYflx
T9QbkpVA/mHlAVhakMC77GkjuBs/eVxkXWS+rGQxswsPxVQpMr/t4OMCYCFRTaTtQxEcKkNCQ4l4
c3ACjvCGEEqB41+BhbX5Z50rkM/l39NizTI3BQmkGIlqPcDLGEdmymy07f6Xo9Zx5JPmJlQ4lHHj
n1jg0U//0bMzVqia8DcTlKnKXRh6GMeJWm/klhoYV6Y0UBXF9KJabxMJK4USnQOsMFJXMGm6meIE
3KC++PoIMRdSZVYx/aTbUHPgfCIo/c5owCN7xvmknrwTE1RvpTKtaQHqI/oO4hXv4ZCU1QEqQqNq
OVfWLWVfbKGdUy/MNUFtslZGLJ1bHZlEagjpAidjXPnLp/qs2EVJ2ZXjSPDg+zq0U3v4i704Ys5t
k8vNV3fJ5XT7LuMp8Hxuv6KIJnnoT+yMjk0kAvTAgrhyUV4NbzVkQXhnFI2SkfJh0r4LLw2ydFtL
LT9uZsgoqgWHN1BvccXvox7kgOO2pHoAeWPvMbLmFUoASAEdAfaFj8hNEpoV9ZxB8IRm6OKLCadU
ieQI8NthIh68MLZDPOsYDqV1OvQuo+bcX9JY8O0d6Q40ih+lOJuHfvxxmwXLqp/pXZUVbSv0p+Uz
ooV6sKmvdZES3n85iAaSEGR2j9rESW5bwkKkcanp6DqpNx7BBiFI25O7PeRr35PPCTe4UMY1K7+W
+AfzoCCDSOAykDM+CLNTNgBvRye0bsBJ0XRDF8WtMtqqMq81NT7uNr1QoM8w2iTzvJG/QznezIB5
99DyuwL1VrsOyx8lH95U+LZ/DvMAUrhIerAtS4b8H2w+/GThvqvloTR+jEVs7HRC4i5z1Ac8NCx8
xRmLk6NpJbZ05FYFTpxWdg4UgrjU3TZ6vkVHWtFIOP579JhG+x1GNL4IT10dnC/ga97FK9fxHmi3
NskdTRp8tyjMXmyiGd/KetmNG2a9yaOFiIIg5pIc0EnBqMz9IZm4GXQICGPcqfcScGAn5+DybY6i
lb329IJ/sKJe6LdJFJIy0kePINWQNAPL+C88k1omS0PpsSGzHdDMUUyVhw00IbIxSwn4ZDGhppft
3UzDhD4Kw8t4Ql6jGangPS98GK1LQ1xKLad1OrhWNdWd3cD6Vox4r0OB7Jmg07+0yADeQCZdMAOj
FGVSzLLV023R+rzK8OGanENygigcC/QoXRc4RgryPHv407FfT8gOo3Sf/AwYRJzTEAJC89k4x+dC
IxapTdOK86/yBUSrLN0MyURxKU813FJTqXEkYuG1xBZpS0TCFgjqsfoGtuQQgmqlMqklMVwUw8jB
OKBoRX37WKk4TFV6+8liWyvxftI+XqN7HoZa3CW0UT5EujS4LQEvkxq5EWBsDYjap4ehKzpwXExg
2JAjDDSfs4zEFbF2kuz2zNE9dSm8w5wpJNS6UoBqV5ihAZg9hgKj7U43y2qsatoyNcT0ZWqQraIW
ST9W6vTbx4sftxI3CZcC1EMtuMoq2IUA1218r5bz27g6N55CVO/7G1/S9WAnbt9UsoTNocjDB6pH
nZcBd9EXFHmBowOIP+CTwzs7JXSYr4nKMbnh6tJFs5HlS6HivJ2/cshp6yDEPif6EnGKyJXKTjIW
zn6YelQn32Ui4C7ZK3+/fkBh0O5He+u80beAhMXUNMpqzuMExmOFZZxEBLEOgyR675vuLCslxf8g
IDSGLIZyhpZ4GsgTMnnHlOiUrBWkdLVLUeoEIVfvW2E4pyGXBCNJGP/99USFDiyJxMO70qBLK0e6
ijkYIpPTdZJ6Q73zWD9lIPxvQYUTL37Hoy3lIqAo5q0erxfA0qmDf4D/NgGVGDcMFPNvbq2gknok
Da5Rm9zj5Pzqvbxz018m15x4pLtwOv70JVoniH/4opwTnVcRKY2Yhe3BWGm6OX/ad5ZaoNkSL8XX
JF/e52NAR/u7ve359duJKvy6qZpf+xAxjQ0bw9Pa6JQ0wNMantKQoE8QFvaC9Lwam4QOpGwDlIEC
+UZqvyj0vOFPjXugq/OMCVa4gCLf90VKh1532fRMZn5hKVpHUWaUe3spVl15S/DOUwvvOUCXhmJO
T6NWnLLIf0W57Po8Z/rMzj0ZI5d9E7jTBhre5X//bUXR/gJPKvcLAjIls7c/92JQGni/OUizIQzS
Andw/xPu2RDVb3OxHiWJ1Pakpiv9Eov78ZcmEqaOwjS66Qa1rCGNnHFD01mYPutF1eNTPZT0G4qF
JltLMGKCizUe4sRmh3Ig458WEFUkQGU5JiHBwSDa2uCLrIii/s7eXkZ7Gp/IzUOQKS6VZmWV/5Fp
Okw5mYVzic/neAziUk0HsVgex4z2jWOwc5Akv4f1IdSyv8+bwOTR0sgY/YEl+5aKI6M5KBsf/H+c
viMEVrGEjdvNt30ISlmRPwN2BjsYy3o3FqE/rrq3sHw2VkhVndYVx8lW1OSeyR+AxMzSPWeyIYsV
4EVfHHptMtc1KHSs98q04I0MIgkDeALH+1Io+3zHITQJm43ggqb286NA0wQbYKifURusVtHQqs1H
O6AhBHCXY6Uxh4vIDwNK6mblcYUlxxnFOoyrp3nezV3H6VhXtemvDndcfJbs2kOv+QDEsyj9EM3b
fItpauJDzFbJboGpoHF9kLrHOcUR68fuCGO+S8oZa1dAhPNcHZuodu71qJtK+TUlP8Jx59visqh9
VVW0PUFHQ2rpjB7j/swu9iAHsyZyENo2WmJRNc71+mnAj0YXz+wPlczZeUS8xVUIISgTHqbpxTmp
cecjGeq3XvE4G1UZHlVwtyf7syscLe0oYK5UfUgbAMymV1G03kP7gm6h5EYL+RAvN/CzWOigKLWX
zembxLciYRfIReiIOgrYf/SIgpZBxtGL60mvDUw1SZk/q65ngUoYMvAAPm0UQxhQST3CZzSiiiws
YqNZKLbI6UIOp/k7P8Ttk6MBSNm0+9mDO/IGWJoYsRoGNs35kQjhmqEL5XS6C6Gxv09AHjfwtQhW
cvjLIUVc0ti/91l4Cy0/eiJP8dNs3wBFOqKO5FrvRps22GM1HitWpr0g9rBtxneMn+PT0/J3uthW
uouRiiT6topHdBUCMowEhNOJXmBNtiEk9meE5WvFhiqtKRmEZ1lrRqwFMwdZxTUYvKgoBPGR1JjP
qsXsH8LHml4SXuZHbQfPf7GOZ/q7SSIAHImOTp+504XdXslQNyH8zP2j8dgHNB49KWAosEC2HfQt
+wAlO/lye4SsiPO1uEele6kRFSwHMb9FX7APLhdYcftqM1gA+FqvptHztOkmnQTZPH0bTgngW9DW
eRSEhGvDpSmRmBTA1sUu4EtUdrR84aRRBtDxl7l+iY5rZDhbp197uP0+xP49ejOghJWBmwwvBflb
DKn8h4bmmKPc6XARF7Rp6xgz1etfHXOyDWgKiz5Ng/MAAa1+kRsZuGrphucp74ttLdDF/AQm2Zct
3lYm3LK4VHoIeV7gKp2hKZODbNmRRIR16nx7/zk/8IeArrt4Ty6xjJap06+53Zfh8hvsLFjeWj1I
NMs/Vv4ep83kZT0xCr9dbEW+n4RmHUg8XnKQq6objmuLTyerz8UAx40B/kdXevuY2b7SlC+6AyEM
pHlLPoar35m4GkbGin1hXSqLedxpniQYC3ZzANiyCmyCdcBsJQGJcwBYI4WTbLOo+y97fWbS8/vD
v7VbIkFi9eOaokjAYdLg00ZzmtpIVuir3DVaZ5ALGGkUb1W+eRjiBP77ULDGTPqPRWPeeElZVLFe
JcfooCvOpElopR29WPa86EcxdjomK/UhcmwMZz0Fd2GTrqKf/q3AyKf71TTh+8nrAcsPkN7jXwBj
LcIYjHwQ0AONWv5wv4QvwhBnxXv2sTY7hdGjM1f1fIhK/3wWabHGZfTje+xjP85oVN2PfkzmPuGO
tbt+UrOQKltfxnwuFKldRoTN2Kmw0ytli1Vwy2EdVsIblkJf5yk2fTfawMKj4FhwxaTwn7MZUMQx
D6swLGRD5Dhdx0Dm4MRJahWS0WNwtViwWrf7/ryciu84+xNyRWNWxWwHTftXkBS6ZsEj4+oRlX1d
L/QRHQERjtuC+qMUMBEqI4M4PijwS9c0T7fyJKKtgiRubbpsDWZr1uWYnX7JbIlwVN1uE2i4Li4F
C5akssICaZfquRQ1Nrerll4FUPSSv+xbH5/k8RPHQT9AebIGGr4VkbBoaBUTq5dzy/rwpaqvkhYI
jHhhGFp31MMmw57ivAWXVtRfaZxzliXNnqtwR8JmTLBcyLUmvoK1eIxtsGFS63M9e3MmDOO3xTuY
e1tfp1nKoS9IZJ8NHb7V1xPmK3xf1rbanPMUL4cGTZ2R497NZ6mEzF/0yNPdR+dB+nx6KLzEFsm5
ZtQxID1LDus5uqsh3waESirX7XyfYmjMfJJb3PxjOYoEvMCe/YT/ZrF8rkC1HfeJgi2a2LwjKV72
i8nJVbzMZkiE/T5Q8bcgQxr34vvBSpZLBVSv7qKGyTDGrNg9bT/8rHCgCqrHzoeNSWRNXPweYEGC
z51k6xMhBUJUSNr+0DJ3AryQoaI63TobN93tkKMLZzAwud5Te1cPBgle/IXu1Rb3Re8qZTuaiYxm
eyb5r/kZIz5GI+p3IJE/Nw+Nr3waMr3k17NEyGRoNYKJoE1atDhznYP5gWwUAbsZPR74vzjSlsWh
wOF6wWnk0g5dewhvpN3DVxFyBIein/ePM9NNFP3SjEW2jhWSso7gAou9mUlZL68eZzbRPR2acNZZ
HgAybvzvxHiSFbhBvqKr1C9rjEK7d46XpTWueGyH/nvMsyIPorXJzoGdbsDlBKoO+nTN/IJIKJnb
hFsitwiNN9FWsxb+k4UTi9X17VDozzTfd5Dk9ClD0pxlhA3NOxlYcgamOcws0Xr6uCdei2EbNVnr
YHMGY4Dxr39Da9zqbHDdqrR3TdTreYZQRr2bedMggIeDEtwFi4U9eW5+SR+H5od+31Z/Gdd78xRv
u5mugvKXSTf2TetgknRgomYe/ii7dE6nIadFmB1v8TMDWybn+gWRitxBpvQdvY/ViysKWUEEOP8C
7dbA9BwRyGjVhvVn5FIKt+BuryNFCzNmUZG2AWJuDUhtXH25gvHbyqxBmY3On6x5p9TZOPSElCzc
Jua8jPwn8riWVfTYYl+pR9TrgkcXYFUs5saO/deSpXTUflya3Irt3I9iOtekG9RkQi71xcYGA5Vu
Zh0fvS2UTRwhYomSehquh5qVO07az1Jhx4r5UnEWg07NYuyGsMs6FxPLEFWM1aHj0hf7NpiSUEWo
c3EXbYedyO5Ptk9UD1PMjYsURLmqA1VhiNlG5yhUwavTzZgHQa9a5iPVU97aVsFw3zB5WxPAlI83
p4s6gmrmpsqE39bJq4nPSGGdP11G7IB8QGNluMS4qyJktEqMp73dM5rE3lOR9LOd4ra9rfHNqVUi
CB5L9ogSN2FjdoexAA1aD3PlCqWuBpt12NXr3UFQFMSxLC6na9Je/CcoebnM3QwBg6tKEwWNpiYT
p5Xxai1qsRRtHa3mVg8xdGzJgcCKk46uQWu+zOHtyTbsBQqhka/7VXBC75EUyaOMeLhozYAoivOP
C2NCWKFagepHnKDLKHBSwASFKsFTJlzULezA9WwVPYGXpcJTcB+opSZwF9dRszPv9ZVBeWA33gQ9
IvjL45tEtXQDUup2jfAxjUNk3pWkFeAzhyM/ZOFTimXWozB9qkyhOiB02HbAbCZthCBkyEYRe0kL
Uowf5Y+LbBie7AglqW0czt5EtBMFJNP+UZzAMNtQIUBVsCYbrPnKVoUuqQ2LcpvfCFnKSZIHoAyZ
wFOKH4sYi/2wCWvp2TcXuzn9Lf/08ilHeuSfiU6TlRAGE/v4p2WFVoH2tdjy7ITQ3VEFYgwcbkO4
YSueDiJ6X1TfD2aO2gEF8zltN0zaOHosfecUN//CcOF/ZVXOIr4d6yUmeRD7FEkILoyEnUpUOPSX
jRVDxX7A0Y5UdeLT0PpQ1zgimmBVodnYL6npfv3SB0UVVU/LZjDoP+zKmodK65Xosd6OUlnWEnT2
ruJENe9Dhqhq8WfaV3V0wSVRKH1X0O3GfQ3TViQXABomSDZwbGCdi4ja/r9tgnwfH6+LjyWpDvdg
nCS83XtFqZ3TjiqwyjGw8RjJ3uLcypXw57nOJ7cpbes5p9X7vx43T2cifN+0CZuvGESujgtFBkiJ
CzOi6aT5PB2t2nnvdBl2wxR2/o3UtV9e2Lmq8bY+Fuk6Z1p/eIlqB0Da2bmw8uw1Nzgec+cGjx0I
HD075cAR2DpyrF7RKz46YkxXlk2vSowh7C07sQi7aeuzpQwmOvu4+aG8ZlyLvMxQkilNPiT4FgRS
a2MHluIrbbVAH9JJffwoP5KBiMbnisgAjlzRp13jlgu+qCVU55R21xuN4u1HIqGa5eLw8nPEX4ex
hMLDUB/kO/k8KuCdOyqJERgRKhMXpO/GWBzZ0ZDv/oqaXaXB+1fmKUbVsRmCHJESLOjWivI7ASOz
KuFDSLaBqug0m/B0o/ywR70xMjn+Z6eSCyOQL4TVbw+wXRdZ/zAXZszCfaaBOcY/nQTZGqMK55FY
2z1ECruTsFkxtznR490FtVbNobnoT0X5evQYBp5ROCG5MOHg5EeNgknFuuR9ZKEPhWhnZ0WPDBtt
9Q+mQrmLNuRrLo18WZHRtGZPs3GwqxjMvzFW/WYn0BSTTcloFwmlO3zXSyrd75mkoORZZOWxSev9
esvn/HE2Iby87LNuOIaBI/Vl5iu8vgeocydM4zKA5aO4POfPCKLVQpZD5a2fAiR4r3/XzwNoLNE3
D2I4PHnA987jil6MragKcYDKg9IGzLvy7S1UhYuJHx4NOYsAxWSeLg208cE3uKW9q5oaqNYB6+qY
2gRdkt424CjWRqeCP7ozlzjzMfq4BVJcYWJB4UgK80T71EUk9AObgog0MFjy6o2RJIQAV5jYuIKS
lLEh3/lx+TVPkogV7Lvds2Qi9ktdjJEOdMcfqCGNDVjxkDZZByGfKRI7p0F2/N5HRCRgzNafC5hL
aI7tY6Lrejx4rS892nQhGN3qq0BboTqNTASjzLaAaUbz/s+w2mxoqhzsZqyDQe+NGKrJxhZLBh2T
dcnSpg0RB+h8TWDR419xk10MF+pw/7h6vmfcDujqW/gpYc/yiccLb5ROoF5v/BAdJfyEfcYMtecx
UQeyEINod82IbvKEojLKvW1dV0DVwGT2yT4BjIHfknXxUfWXlZf5jDIoXsVtjqxVtaH7bMPq5xFX
z9uZ32ZVem0QiQAVgGI6WTaJtDRW4yDyK9fClqnA1ocHScGyWmJQ214RD1J8sUlwhuSdF0o+mIp+
3pV4LoN3yumhJQBeA1RuumYGdhYmYOeiCcF86u6stYvCeLQRlVMDZbzmePLs7bIWePx4qP5L50d3
3xH5+uXk2JO4K+9SBdDdS7Rm8PMwAQrKE3fKrjJKH95E1GJO+YX3FX/TWT/ta+Ms04T4ZKjZBIn9
UtfT6iYiDeYykdvJfTf0TAYxrwYZMnrjWPIhNEq3MqCOzbdsA11zxSKAIxlXm797w9Z2ToV6vNXQ
p+P8zfpv+sF3ZoskjEUuZ2yjJ6WyVQthqD2wzzcu7KgXVpDfYA/BsHNBRqqIPlulMa0TaKYvMHEQ
wrIPfJvrfUvIBdHy8l2iHB32lC5VMs60Q5/V6CVk1IBOcCAsrFD542mzuNWRFrhhk6XDvT/2VXZa
khGrkEUiZmR1YSV5UoiPYB2N/4UaoTdYJOUCbG0XompUQojZLt3C2EdohlMEXCVQXjE12NhoF46t
Kv6hmrXX3P1eRkDhffhRQYndd481fiMOGe1guy3GUV8JYWttyDj0FovyTSUHhUhT63b+HxnXMZxQ
mMsQ4lSBQInW2t+0VAsGyJ6aPKuslH+UvmC/BgJ+MtcbF5iyEDSSLXBZBacwCaOLJEPUu3726/ie
fpT5eJOPa8wSyxZzJHCVTVaiLE0QLxGpHsvgvXDOhhva50+TcOKJzTuwcg0R4G+lJabd1bRT4bIo
ryTGltZ7r4crEwuXtkOIZXqvHgoAx3aDzKeuFfoddecPtnmi5MPBqlbYOIJHSByOPm7DdyWHyEbN
obr8xp/wbpc/5hrRo12UDsn/RmK1x1ur8lzl283q9HYqZZ0tRmiyvxrjnjOLV4PcsJ3CME4HcgJJ
AZMoT7rOW+vgSVZKMlouFd5zi5qfoCEmc69wbpzdKVGJzPs+b1ILjFwXR/iGyDNp49UkZpVY1mEM
SEiu0u6IcO5sg6koGlUX9Zvc8vG5d6yF5XsMzKzND+5lwMw/4SqlRUbfU9la0UvT9QLa8m2hYBvc
HtypSmGXuuTPgbGeqm8NO1kpauGxLRjozkEqwi2ghLA4S7uJjzIllFtDbSLV6Vls2Y94F4PaKHtR
8EZyuUnjzvYvJGHnhdAtswhuBEyRZbFqGJ8TUB8waCBIzH6fs0iKNtrufl15zfWfShjCPm3RqexH
1gZFvN4r9w48zoH2OE1HuOyMmeIvvhmPzYRVF9T8QD6Bv67Ou1hqb2oKKwWU6Ew5tphwbO9G8GNH
SxqshRlfQaPerKnMq45ZkFVEb/7mvwoeTUQHOYWhMzxQhw0Q/66ZYnu6LRV5xnLlavl6vXzco89s
gQiUAVIplFhGHG5fbCFSdrv8Z0vuOptSytnCz+499c4goddR1TICQh0g5a7U5gn3GIDva5CwtxcJ
vlAvS7/khnf98HUlXEBcSdY0SGQMzSB3vETRhEJoaPo+MkT2839Jc2tK0+Mc34a8VWfkEw0xJoCG
t3M/PtIFt+C1j1FUsl8l1BHUW6dd/7rUWhGoDjr+GsoaWh4FSDADAm6LrYcMuJi1IOc8RXqKo387
nLNPJsVMlBbpI9+SeOpwo17Qbe26niiLdUZxzwLahTrfTuxIkvR6tawznrBIgwfsG+bRF9/lAW3O
4eiSB1zpL3G5h3lcv+xLBpfOWDblWEsb+LebuJp4lPPf9Hg44KoiZ53soWO73DWWak7D8cr5c3Nr
yLWA7SlMyaSkYIbETPIcjLsGJjEHgmgSOr1yXL2ZLSn4D0au/Mlt9WCTaBE6fOc0+SGAqVgkZ24T
gGoJZ1dcoTLfad6YG4nqM3WjxAZ8XVgMzNEYv4AT0IJeDtZISIYsF67P4fNAh5Z5mghGuY8tTG6x
fR8C10RyPfTD4LiQ3C7NFHGTH0VFsUSwohg9sDgxVNZ/r9hSRtFkLE+KAXh8U6ctMgFLghyib/1m
2NGSj4pY2I3CStL73IGdiI7lW8FWxXGs6LetL50sFQ+icyl2IiHNPDRErwSoWOlkw3XFMAboal2v
2c8SrY892c1oV4ytIVQloQp5j1aAK/pdIj7qdNy25hRYom28esemr3BVUUgWZ4f2B+tcerH7AL1o
zzSZriLP5FIwHZnYkl7OdCTJwvf6chaHqQp2FXv4KBDq6YzgzLX+CIaRqg7HSRPkaw+TsXtbtW02
Jh9fRWnvzp4eQ8VYcfHO2b8Zzg02F4fPQWoU8lK1Z7zG2rSkYq8HJvKkb6O0FiPRpnqVtNaTKI9F
j1Y/VzAB9rjK1zG0wCc0hubkh3lXmx8/cYHcidjmQNB8iO6ngANhJ1JgzOqwjF/mBNL/l7uQU/Zw
/4owD7sfuu1b0RaVFQN+dWnxqsvfQx5S2mDMeqa9XLBgsgVZNWFqwoGZo42dAtZNSyp3e1tb5jlc
Wj6M09KNgcrnqFG5tNhadHguis/mXWU+4+I3nYiyeNhWX1lthZRnupz32jKzCyEz2ncbJs8K1yJ2
LGhu18bH2sMyBLH7J47+lKDMVFbB3Ga2YxO6KU8vKBybDhwAlnzhE20RrIpUQzbhKyJU02OhT7Am
uhtt1rSUwdqzBlAxPjSYRfE9/+Mpibmr6yQT2Czv3fGBvKR0jgmSA9/FuqU135R6HeAL88dY1pRQ
h1lzdL7JdXO2DPKbnuTuGuBDDRIRGzSpoUBs93TRiwfjC4ab1+WeNVkV/ROhVbV9slQjk/N/nEua
EzojOI+lzkqbshrB+UQ1XL3A/ARslUtyr4DqC1WG+Xh7eI9qlOnGmv23vNjPPRPQ9Myj1/k1H0AS
qKGeFjjlLLwzKZ+Kd6bA26AQQiNQ3O5FTZ3p2aJD4swj+ZsPWoSCg2kYW7lSj/t+LBJrDJOXTEc5
s2Q5I/Aojm2EWr8RgbkxagwQS67ijC9rs8oEy/HBcqeR8njIy9YX3TvczT8Vjxll8MI7XrFuuaCJ
xZ6Dmhiw9eML3qgSiex/U9YLUkmYxJ/UOdINCT9E1Pahte5SP80vd7jr2mlw5/plkZJmYo0rQ81O
fO4zsp1SP2R24CKTXuRWVJco4iwToQW3xKYWQ4K2QeuDaBTyRRjsEIeHFpoNxKdsIVQOuyW6SuHh
fp1FYXokoMLuuq58a13IizOgi+EN/ME5KVgRaxONW672453npzjYDSrbg8o0xRQSdMSfreh5F1+0
Y1Kzfn68f5rSLSUjRUURfPXnCBzkaf2rdZB9AjgJbknMGcSCJpNgqLesOr/H+VbXGxOF2Sp9i6G6
rL/y0CSZdPvzDdjlA9DLf+epOsgb8Fdw6cEYLPb50FuA5mKl9rGp+bKpxc1m2+2MGddM2wC7Rjw3
53P6nzjgBiQAcewiLki/l3aGoe+5ZFgmmz1KZFYOMhL/zGCDyk7wxsh5/ygt1vtwTve6pKqG0j1i
h+B95b0571YH1OI45cZF2rWM0g8O9Sq2Q9aDLwsHBajce0Eo8azuUK48wRtCdwWzALOJop0pf/Fa
ov8kvA+wWxOoXRzllGTGD39dLFZ2LO9DkDEb739GhqHuk7RDLbqazPDCAL7lbEoAcoThTdW/jFjF
13Wylhacy5z/qdaNjL0vDIS0wdx2TpQTXHAAj44HIHuGoWZRlpmxZ1KrNIOgT8R96kR0QbV+FA9X
AuvMRoVsSUE1Y6bXWr5kJmhsz8CglNCNLvFj0/4TN/iJeaYKzNFKoYn83yajxvitVBXzHWCxVVUe
T7MagZkNbz/xBuc+rT1wBUu4xMpN+lHPskDrP7ngj9T+A9USRt+cvPYiUEabh48x4UoUzmL2/myZ
CKcjvtJhGgyzhFceuAzwvdM6Tahrqspmica8QzacIN9cDvzr68nil5KOcETjRC5h6uBhSsXLRyyK
4K1UCf6AHsE9ic2kZ/7kTykMdJADBTcN/+Bo1uzxZ2LbnWYq0rY6yRYUJZCB5O+1v2QcJEMBd6OX
FQhkYz5csX2nonR9rbU6XpxytKFs6ioSevZPKKdQ8DeYqvfg8b+PptLekLkeP0MX6WPHngWsBFlo
6sI7DHANYXNwdWEEgLBmItybl9ScdPp9i3NUo7H7E3eKQ+GPuum/KRFzHVWy1v1MMTxRJShwM9FH
x4qdyAHDihuwkb+ZGIe1+fMANdMeZrUShzZ2KVewpFrnho94baBy2wrwncbYgSiMEXhyZcUqUDqZ
/LxNAI+G5OVWpZWLeYA38zRBiK/9F51toDfDCZlBwpHmKrviDsLrIBNEz9UxIL5O+kbahMElJqXa
vW9wpHi+2fPQL8XPvHiPlsqWsppPXHCPX9l7uTgUU7DT00HIBeQlJ+9VQ5jbaZyoyg0aLo4gnjtg
TdnIPAcxoJ8LDNZO87+K/HmYd3jc6tUiy6EDAuaCM6QavUO3oBfBOmeTR/OmgrgmbQOHFsK7gwa9
lyoGBkpLQ/n1gnnfdn5Je8dxH3bvx+yZz4koaJdYj0pjg7/a6jyWlafaJVyzLMfhF5MDS/Ka04m1
w2xilkHatyvvSbghBIs72ZPbSXBBHvxlsmJrYguwLlsTnUyoykyFjOnzpaAIdgl8o1LaOAq37jO/
bEBj8+xuPGy5iSR3//wZidLEPbz8uxFaYT05JlknJ1E9N8njG+HsnExsRs57vcfj0jJ/BcsjEldo
OSAafSksAH+LkHYCzeXsXNcWVW/s+w5kQNZNtbzksX/kz4IAOCO1g8itUg+NwCYf7u6on/A8lruk
O7yrFmz7I4+GvyyibdppHAPax2vYO6lER1n5sDmrKoQV08G7Mk9Q+3gOb4uXuK26dtWa+Fk6kcqv
Rx7JDZwE3IcFXhZduKiVhXbABSyUCgyrqlKAcyTqlyBVlKUwwJ0RBSh7sXhXMRagmGk3rvXBwNRJ
3ZhdAD0Uxeu92ZYHiY7Xtj0cdgU7d9YxSqAeI8xnNILl6NdN9VHs172oirDycWEU6CNOtqBTMBF7
h/sD6O/uI663117nKyxqWwOHGxzbN+IwRNM4wmdU2QxBK9LJE9bED+9OA/+I90LawgrtF63r/q1G
RIvyhunDxtXVlqvCzwrNzha+MxaRyMErpxhzgSfabj4w386R9e0XlbxtoONsivbhEJHYie98GtGr
G6NsW44YEWsMAcdqEWkDQ6hPtnRAKJJvTCp8TCZYz4xcn4fzLttdMS++TYjRwE/dEnJEs7O9xfO1
znN+XE1nhYnOVYTUnRA6PzMDy5KRi8vfUQXJ6801LmCjiIyHQ3Ma9/1PF3thiJOfBeWbKftWxl5v
XxXPm9xEQcV8M1hUltIjbdSoWuTGYIWGo9AXXY8tCjW2VJmm0uLy/U0iOjWdAidWUL1XMAfN6V1+
C0n+/I4NNPWHZZuumjCmN1kJ+NLHTWOeIrcSyf9pl/URbVUyJlHQOmKyKnVLqvzl3qpUE0Weezcg
nWdu22pM26ydT8gx8u8BgBnu+fRr5vONqDUtAz4YsUnHHb353pE8Ew3OcYvoulYgA1SgxlOqeHo6
LYIva73amYUh8nTts1asEZ+B11DNwbEp47yLpZSh4wFrMmoQGZeGMGcFduVbC1pBaUiboIRz7tGe
5gR/U9o3P7fTiIlcVAPlUHMZxOGni2vcdwcpvO3+1OpoTPdMaE48JfM19krSU7jRDeyBAoIfQCSW
oudQzc+tPHHQQO0d0cAu7jdn6K45NjSWvdjgvY6/hZ1UGVy3wrYpkJvhmxmL0osX9oqT2hQLVzOq
u3xVx6bhfVz1gJXzylkW1V42xs3hbfZb2gHkPi8/f71k8IkSWfXIQZQ7V7Su6LdRWu+jDvyuTPiC
G/P6PqVO5ryA6sJ2M3iBDTzb+eGDrB6QJS81RkLmRrjoUFzqJchNm1i8bcwIKsDEQP7QmD8bsayG
4uL2IBa0iVbKZh40dd+0BIPF+z8d3D02jPNX8YgMn+/joqTFREXpw160J+ZU4eU/oQA3HUcfGExu
gLVPPGIdLDY+Qc2E2n5Dtu4P1yGxdWiVQ0s6gClLCYMstnc1WW8JE80Pk8+8YUDNHCOdHOlL6S0h
Z5SBpo83hudNgcS4mCjjk+1ekNv1q9XRT1Lmfrs2dzVZtNpanhquFespJbuw3ZIP8x+ycprjgA2m
JonPJctdYjXBi77enESYc7wjNfPyJOXsa21q8AU6pFnk0y488loZ2wZ/4a23lT3chK8slAo//FaF
gl5+KPjIYx6UW638XGANlwZgBGUUEmFObqs/IQ7NI32FczCbpMor+P0i1KHCHInmSR1Bd6JwyivG
PZxTMITu5mkbMyvGT6sWBgghEVsQnEO+vFPPqE4D9V6jS97jSMW2iDKgOylt8LY58wViQQxHQWld
vSesmi3MbeHpUnAKgqkOoBeFNQTb+qxUXe+Tw/bsZ6ysGuPD/a5dREZkpn+VxVqMUUmf1QkjaU0f
G6u+9Htug9T5jG/WYGPP0ADEhr9hd3cuSVzeD0/z0TtqY7eXTd0CIR+m+PolIqOXLE8GEGzZ/xJa
Dm/VcPKNCtnUL34Qhccv/j7tXf2HY1fZvkUsxQORUxf0E1VQ0dCbdnq9zD/dpEOO20j9pRDN3lfU
Qvr56PzxXDQ/QrmV/aPpa7YxKj0dpYNwBqQqUPjaqpXn45JbYAgzAUmHWYHqWJ1DdfoV/9wpVqox
u9/6z6KJM2pznSREtXrHcojgJlrR4OEpaZH9ZPzLmkFqhPidn/nd3kPwx0jqWq2iglT/b2n+F7g+
PagT11FtqESSxJ0KNKF+DxYr7ivzRosv1KsC85fLe0QvR/plRhA3cClqsJen7Fo/lieOGPWHwiCO
oNBq4P6TOLXQAkBldUtlfuFz6B93pR96gd1zZx8EyvnfDUnrhxJ1AUw2rPXrg7ZOwbsL5P5HWLb7
IxJRsW7HCtaqa2s74v6eXLt0o6tzv9FBlgiaJvzbPonWfcHdCWGNbQ28kcAXRUtj1U+5fp03cvmC
wd2yea1FnfOKDc+L6MnSybJSfeDHtXmVsZuJowIGCQ5WxqX2EFw7FOzLoAcIwTQGdRCBzuYCeSuJ
wcHod+dUQ16W136fFKY7OdEkPvJ36l7jxUa7foZfvOCQBlVEVVLwmQBPTVeKI8NaA9X8SAlOP4eJ
cJ5mJpvAGQNEQPwubXkBNmBXVBecqdIpN761LSRhnCmureTqffmRiTdnABpLCsy/VK9vJT+9J6Vw
Jq0Gu8zGufwSTtiy41Z8g6oAMq8/FKEXddmGs8v7LHN6icPqlYuVa62EC3Bupm2XjUlNOj0elRKy
XidBQIT0rLdWyB0By1OSoJUso/vQ37JHkVjLKJC2VUn64d1MjdBPKNYUkS59bMbo6QkrIv1maw0q
jyD0P1SOlldISLyw/33ERxc0r69dXMIQvQZ3ZNkofWwOvFAxQNSNV3XmiIx1NN+ktWNwAtcATqUH
BDTs2ZhT9zr8EeoM78aJuEfeaxedWsVjUg0bvuiXSduYfUiXcWSf6nJtlHwXEKPyDYEg7HSofYfR
Tuq1AxDzc884z6P0wGyz8ozLygQAuiTurcSx5+BwlsDaSgJD5JT4eh1N+SAseg00el0CrqkfRDtA
V+wIPoml/1MFaa5IC1mw3/pXc+7O/iJCZGsap0q/Jn800TV9HAwZrXtGra8FHkjfs2w8BzyiS7sN
baTFHodCuaTh0eVeBjUzi0GkAJkLwN671h7J6JpWeNIsLyJ58Y6FLOvmgXtPPqklhDVPb1WJuiXq
XMGN+6TmHhjF3WZI/oW5SQRLCvgoZ+S39ttV0BcVmHyxKGIKloI3hrw3YhBpnYqyBNMm7g7qeosh
mu4m+JSqeLMX3TGjDNqBllogp3ZofFGIz6k+8VQOnxF42FPWwzE7/ttuY1svNNvf8K7bghoha8G3
Od0mMfUg9B+Y7Srf4x4uGDiCVIy/Ebvq5wpkNcZLARlBX4FyFWaW/7+gQaSBFglG1ltWqt/i+bwZ
lQjwadLT825g+BLhqgtZdLJab9M4qGPbCaPGfF/oEz4xU2OgHu2D5c21Z7jzUWi32/9lmBafB7Yq
TpNgchF4HQLjukkOOZTE3EC56yWA2W4YvU2GTtVXXW2IdXS0vRfhON12fwxIzVwlsT/GsV5e7hf9
QYXZtaOEQSxXNcP4YZQvDt1umn+/Q2P4y8QyCz5UFZuTG2vSFU9yuZcPmqNzSlzb12FUN8d+QBwQ
bZYgn8cN8/xLoOZVe0HGFFMfdkNYLYM9BEkvJQonidq0E9SZZn49bkVv4vjZGeoaavl8UvXeatqu
Nnp2GdZitrIZ/b7+yeSJrPBmCDZIocTKNFY+L2r3tKSWUP6bc7XOeQjOs9MmD52c3kknJksougyr
EugfIn9wYNQGdsMExQrRMGu+ZaTXJacXOrRdS1RL0rGJUg08n6jThbRi6MQ0a+hbVs6dDSq25tEI
SQlHpiVuQt2fpR0NOihF3ckmv6pnLA0QUiMVK+xoRcSHTsb+6ER05tgufqFXhpFJsoDdvrcwURze
02slCQQ5DUdFpODH7ihUIt4pK1n8DuaQz7wTXMxRC8Otfa9d6b/4SzdLaYF3CG8TIJMzIxVE9Ao+
ZBYOpqsyHVIrpaEm/dR5HBW5/+OwWg4++8Gv5sH0WTlMpLQgizrCTS0lo7KiKVrtSFv/q6Bgfk6B
DjUAz+eWV1IwzEC+eNqK9vgZabvGWvpsNfLUdMBfCdS0bRfi1EychCM8R/0mCkWlt9DFeywQWm2g
CW68c4f2TwSZOOMCRRxCdnvNBSkVbsYEpmTUSuuOA21bDtRQ2wiFfBXJmGNze2vbYkswl/XvJVig
VPDQHnCF6zl+bC92TuSn+s7TlHemNa9jWQKHG7R6PnzGrRhCyhdANbUrCSHSzOWE7wGLKJjr5aTw
gNq4pu88TydkepKEuMC83wILKf5wd669TSH9+EgdRnYD+fQSMVAXbkw3ioqfdFc246mMO85EQHsr
QA9e7DR+RP9wGnFUX8ceiyp38mW7J3U80FJ7SHVokoqHNGH4NMuRKHa5JdaXj3xQdoLc1R7K+1dC
eE/t7LLHWJklDUMcV9FB9MlTI2DtW/Ooxc/B6O6tzPqiywJE7y4Ppoj/2AJEuYYCRCZFDK0fo62+
1at1kdrn74oypzxZmXm/rU+DFVxCGWeefIn7k2kZ0F5+94SpAsN8LbLY9YVCcunzEYFNpipn51/u
Zk+WSavnBcXlHumoR+RlDCIKSyzkVzMk4ezK17SwnYQUV3/jI1M57NtZo8zEPXdEExwHTULPvUUg
G0nzo23hrJvPfdW679X1YT6X6y5baLy85KQy7QFOdRNMVp2E+hBJrop3d1cbLCml3YC3WMiNPQRu
RSjaEHiP2EgV0QBYvjp2u2gbgQmq3BDmTL4Nwun3HxtGCh+DoMFxRqL15+Pf9VH3Ke7awYujIKkA
Kbw0pARsRXMfzCwmVX/Gj1hBHENypVC65vAm2EwHoJVqj2U0Ao1tvThz+rd+6BDq6DSgvCddZ7Z3
Q5W9WTeQiandManHQ+KHrXm5KCz0ONhPGmzbQ43+dISU5Vqvqui4BqkFeXqAVMH1FsiRKPB4vTGu
l3c0c4QBlt1Rzeo0DX0RM6euL0VTggShL4OiseNjU/wr27JM85cmmUpp7xxTuu2rwhhJE29z2V/m
8kXtZ5SDErXiU0V5l8eISTfGL3IZsN0YJhC6eWK1Jd7pf0HT9DfLoVFefWxzMPbGhW0xRhr2H/92
Abx30q5219x3HEVoCplqc1aoX1XvH62C7MU8eLwscISu2SX49fdKVex0eb22NCggNo9cKDz5+OYL
RyGJG1JaIh88QV442og93pqJSbP2GsQXp7BYJN2CbzZxjgrTLGTTuRHyP1yXR0y8ew27Ab1HPbmJ
0BuLBwzjwUX+6qBlL2Spd4uIc4JLdIVZfBmqaPlzqG26bLzEhwIW6mefUKZDQuVaxHEHs5ZLjRTA
NKdmjEEHAQsPHOo/FH80RP53fw4aHeU+dmx3TdcNsYAfClsXrKlFQlDXuRNhsqvn9aaDo/zWqFLn
eZMfhzlteALsIBPDqPG77FXTAkhxd85i4nAnm8ecuoTltD2AqkZFk3r2HjirD/m7yFOKoZmI88k7
GxjKhFOITcygf0Pz+qZYe/BTcIO0+nF7iTVrR7qPsm8fKg4wwa92dehFnN6Glr1c6rw9ppo34lfe
W32sS2ykTR7Hoyqux//9N9inBXCw6Lll5AVUm9Cbhe3wuiSRZJl3A4gsdK2eHXkudkoCrPUD1uf1
aKoi66Ps5Svyt9+uKceEitQeXGZzNYWIeAZndlXsWSdDjateU3k82BH7LmfFAcErm2OdFe5HLGcT
SifHavZcoOuLJ3DwQWBiaF++PZtPgJSSPfyGi3TqU4dZvtOzJxLUofsd9dCMw4Apnd+3TXofbXNy
KNO6An9c5Zx/OqsZz/H81vYAkCeK7iVxNgRShHDNfOYYFXiCQL0A33zt4pBfCrbpbXBbuWRdvz4g
5ECgm0xYWM5zTCNGFOQEPXNjSldcTuZeXq3YNUumbimIjMIdbveJPGJJL2e8r9DqL1uvz9bd5FB5
q9wLYYloDTeMHNgXiA5ucjiGRJPw2zallyC/+jAiIFhjvFsi0GEdm+/sIe9qJi9We6KRTwI5uYM8
vxf1YemIfTK0J/aSReUqOonYB4rnYyWx49JurOtGlYlk9NIkjHWudHs8PnNWvV5txdWZnR6qIXdA
dMymrXeyPnjK2dBuI9+z3Y+k1gOtxZVVvYdrlPgDvj7k6RyctrZOa56Ww+k24oDpA1369FeEr+N0
WWPvH9S7LXuvi1ZuZyPY61llYFnDLKEExarF+TXqrrmalVQrYEY9Ab3o32ObkPmH9t0mppuo45Wx
eZMV1Ev5hvE0K43SUlaRSz3DepHHyWiT/wg6h0byZx2/w8OJU+pJNbuqEu360HFG6mMC1f7L+wOE
wMuAjbDjiT5N8IPSEgg57gDeY+TXJ8DfcouAHq+6yoWpxHJHSP90ks0R5AMvJfrSsgh7g9+xRb6g
WDI+Uox9cW/lZGHGVnvdAHtClTGHo/K68cIH9F4933XjS+nPXYy1efmjl7/itCvr3cOGYtDcHACa
9jBvvaCNbjH2I7K9noVnIcmPmuE//AXPwTy9fxPPA0z/flng+/7HBLHwkrFmCpQh349Rao3Vl8kf
JNq8hv/j3KzidIklxgu2kEkpej1NezE0rTqjnKv1dsMU2TzCvL/ZEPzxwe01ES+5/IfEkrWxYEso
D+YOK/Z3y/HvTAHvBaFxSQIOmuMHzWmYmdQrPxavk/MhAUMG62nzApVmbYMZwRn+5McnkkIAXyDX
4RUotgQ5zaZOqRq9WevmIntq+6c0ANtmi7pH8kOPFUAFCLukLThx7QufV2Gv6Tz8d5/m68IQMLE7
c1jObqsTIZTsYh0qjQzp5Aa8HB4AfCC/VSbJ29Xcb6uQVAxFVJs9BpUjbwZsHhvFrRu2R9PwW9ZC
EoQY17YrZMVS22rhTtaw9mVVpNGTqEGmTxCr5zlOWA2bcoA4EwvKYhZ0VpMk5hmT22+0GtWjb7Yv
HalI0mb3Hg0Glyq3e59C1T+PQyXDiZibqMWFUDB+gwtO/8l+rRpzDS2YnPrSY5dRpBR/ZIjjYVAy
Y0L/jVMMz4VivaEMmkaJmMG8TmgiPzyS1xHJLH7ex3OO8Bw1fJYhGaMUGiVHf27IgNnLDBPQkK1u
qgLgS/+iJJZzgNJf0YZzPc02eLQOh9EEa/662K1TBHieeSE1aXeWHj9ezjjT901CSDNF20iCQH2F
oII+4zE8abMHeJF8HBfGRD2iO6Ohx4A1ic4ZEXzMSmPVcrLppfnspwss44qtgjgO5vMCIxDUp8/h
59iJO8VTtNO303qAa2y8DdldOnJ3ek4aeJHGxmbX5Iaba+SBVlM026/hVO6cqwLSPHkae9WRKHH+
tpBxd5SjitxwnACIttviuPvPrH0wg9j4isnjmx/6R7YqplRQg1GUxAENEJNx39YMVpTHjDQPpEhz
gYM59Ao+uht+WKBVMiOA+h2RumKTFAtprvdPkHYav6MxdLK0y8NSeZ0k3IXeZGOGtxTYC+qp/Ums
ztpK/OaDjEN2IxTf5OI3+kikELsuALmo2RwBmZ1so4O0ke4ZgTYckJEllsCa2DLbWuq6YegYyWJi
mDo7xy+/T9RLUVeAQ0CI7ENHQt3dhpBNmjKeImzmmH4LWykjfeAah/xXT95ltsnhrcJ2MNCcrOCj
CIJRRzYgdTjMrwMXWdpYjX8shcheGwx/95XevWusqJzSpw4XlnuLHISutYcBUbcQv0MxRptfMQPO
fdVFdV5ykM+EMjbi/uF7ckC2FkApb8flHYmw+jF71Pg5SykdxUHxAafu7vPCtrCtlcjJKBaNg2OJ
2rf73as1gjC66SVAG85eEjktk3xBVRpdQDs6nDChHqLmTMK6h/+V/KeW5o/tCoNX2EkNzOeKTh74
uuCuE0/1ORhtsXkf12P7tDbsEJdRzY40RfNIPV9mF57ql2NN3NGAlFXLQUnbc3pWicutHVzpDRQ1
NJy9BW1TwKK0ZAuESKnR85BL6aDNwldF4IkksBWMjqrZL5JzBGGm1wFtrrVbPYSdsj7N/xQPNhkX
5sVf7eS6FzWmJ6juTKvihnlVTPVz0XMdsv2o9S9w/AgrRqW2favPrQFvpkshRh7YICiSz1kpNxqd
HSXISkL/wN8Q0hZat6VlHE48YVb/11eSc+G6soqpeIDbn0UBqdOO/OFhOzaIiQ/zZRbI6qda8Y5H
bciQZ3dEFyvibIoCZlR6M0C0RjN/3h6QqCMyCM9ZxgqZQWdjQi//OLoKXudan6TOpSJDzC0SAbsh
LFJYkfkiFgk5eTYycVRr6M1no+T3WJ8k1yx5HxnnCFAmDLmlEGzTvLHrpcTAc/LKrxbchXsZo5Jo
0ARZUb+aPBLCLPbNvy9CaZsgwVEUceBAmcCZ2ncib3ItZMf/AjUCI4Tkk3hcBPp0IxP4LdpISsas
qrIR7n+9IZPgZOlPQtuayUI01pIIx82mX43c7RstE+agKhNC8saI10TJRMQSVsENtPKap2/e2Ehs
fAxlEYsnAuJib0Kuu+4voWzIrTlgFrNlfQS11Uz9p38XzaQepb5b7NjQ3PGXtUPQAyAj/EpS5JDi
5MPtPXVwiWt9wIQaThygQiI1Sxo+yQNj43yPS5f2eIcyvRy+dY5fVRX6cr2iXGiBBjkWJG3AcOwN
+gvM5ppj6g6zl4lSU8z6IwN23c/uaNXskdlvXSAC/JsQprhNCAoukAwLPhzXBPQZxKH5jOsw0YP1
lMjlqdFMscNg7+cHhtuTZ6NRw5Mz3QgD+6sBDgwsHnQzp/hWGbj43V0IqUEhYs0Wu/ASO5SS2kpN
ln1ng2zJOXp1KC9bKSRN888p07mK8wSEh9AQXdWS5ETU1nd3dk9/gGRpnIaENTCpweoPwd5FrMK7
8GMqqxpKiit8NaPNk1NJt/1WNsEACwzFuSnQKVY/ecqDbH3K+3S+a2KURzGCJFVKp1qIHuj7PY8A
xdb45229ToRp2a3pismD6vcbqM+Po64xGMRscM8vBAcs6R+MAkNp+iqMvd00Un0SA4ZhzZWu4pY+
F+0WEywtOyGXslVPSU/OL3UeEGP7/qpTczGwpKLNkXU1MvpEIxS0nnfl0NTo06Gn0GXapXRuV+1Z
mRphcRDBbk8u8Lnw37AJtcBp+ijmo6necobMXwQi26z604r65T4baNOZj79+nVQg2A//ZzYXGGMB
PG/kQw3lWpcfdHBnkarLyuDWKbqIMfUYBzwVMLSMS+hjfpGRr9zRDYCaIkhxhYT1CtBFic+uFClV
qoWaTJIRueBiRCFv8NCdZhy6dZbJOxH7mAOO0mIc3LM9ZdJ7QwGffv/Zr1HCkTNP5QLnEnMcQfkk
p7QfLxfSLSyygI8tC7SU25kifCYQaphWZAfiqk73fcpdGy0Obufc0KSTlnBXe4Pw+OK+ekGhSrA9
9GphQ8W4SDJOXNz281ZUb4ChBsfBR6qKBpiFKr16PpflxoWersrqPP58b4I/4T7HBrRbteZbgQl7
qpAI+E1q9+Tg5fl3rUG+z4i4Zfhf4pnIU3fkCQnlInEj7tnn4t7Ea5XegUM5Y4tC4k2iIzr2frKw
83QQqBwqMj+uxwuXzYpZFG4okYXLqI0nF9PuL6oSJg5dOXZ5zH/5ryL4wQG/AxymFg7CxHGTm4jN
+jtkrq2R4VfGX23f86v9gL+jcLQ4Kuewf0ekuqWu5bNn1KmlXoIf0ldhCGiQzEzUiBxAQSnsO70e
PmCoVUqo574MduhuCdiGpS9G62ZeL8+JLmjDEwnsEeDgAaBLcaJ8cXpE4PKpW/8GfPohpit5Wngm
okO6uBZnVEFGk7l8gayXWe+hyOAUaaS4r2olipXHqhU2wYn+WBUAZoYiNw7NnPG/tIZRCcWw2vPr
fqHxbsTjaTXs6/zvT72yaF/M2wcYojnxbKXPiGpZksLQn3DaqeaHVEY4p/bwG1u6HcRDCi4xHB8o
/mRaXDYthY/ILUtz4xop7mtgTuEEfs3XqFClMPGqw/i37Y4mfWnlvR7iHkYj9Da6ScLDettaasPI
0x681sWS7ZC5GEuxjXYVB/veGVJ6Bj5rQ5nPSo7pZz9Kxwb8vFCLYShBRntgdrszzaOVPpsn6SAd
Ew04B/gkEHzb1FkZ9LvrbZhprIdoL0nfsGo8vyFzYIW36qci2fN7l5cHCBsGIcsPyje/ddjIMfEC
hN5MyvCrVLc1O4ppF1ugekvs1AKgRz9fYHgM/FMxoAUd714eSoytom0gNntYJtmmgejAQPivIKkb
wLMoSZ5wQWSX1EaCSbj6X+S30p83h9t73gxb+bHsorDForAyTb14q7qYhXLifYb4dT7K8DvkUVxx
K+LIAa5Naa721BSogAMBjUChPhw+CwEohNQNLVG+dwNFZVGJizmy7fHJPnXDSOQZ6+8dhwqxL+D5
Ln1YiFHqMOdWGf8AVt5EDG2wwyNqRUGVaJ9Sf8SmgcrNXpnifHkZosB7LCL4JbsOOKroN5jLD5Fm
M3mu5dthq7eJri6EUfIRVGeM6a0Xug5rieZPsHVYBO0JdZNKqvJMUL8PIBuUxS0aoEPWKshydzgo
tSwO3hqXjhCeWq0VDnJPL/w/MXTVzMQjKWqymdoKCbIRBoRLsjw7QKeQy+OLlwtDNRJhon+1mSVB
lzEP1ZRjl944npakmxVH9sYJZKDClV/8h6pDyPx6ToaWoAdEO442NN4m2xU+ajlV8JqSMor55foe
6TMGRpM4DdbUaBu1kSyi3k24tt/HaXWQeJhD3pagHAT8kC12i5hg1CkhzJHxH8QJJAj8xcrr3lLU
W533vDWEqr2ZDh+DCZPVx7xgOayy+yss4Grns1faTZYGB1Q1JNicHT3BImM/Dq4iMlB43lWxsCt2
b+zHG4Tvz0EoEzd0Uq0IWmCukooOm5OIlqTQ+ZQfuwhgXXOcwn0DDzCgsANTkEWSAAiQEwNqEcyJ
VVfjJJ+UIiW996w7JDK8o1jd/S80utxrXePjGex9KA13z+UzPVzti7i2KMGOxcXjiYnVBTxa3B/W
0WqJS+idHdqoiKWDh6mbW/3EpiN6M2B1tTg/hvPHIFL/DWzZvVd+prrJnvF+IyTdxcJnkficr8af
jeRDbzurgnBUS3kmsTc1aqSeNe2m2HIPj5Uyj+wgSzT2pYdzPV4X1RtfzB/hmuyc4s8ZK60zEn9S
5pZKa0J7/IUTFDK3UkuC6Q217DolSwfrBjRjliEVfC8LAt5dGBUN/Ykp21Kl/XfbvpCBotG1QDhj
WdBf5aVVxt9zzTTmdzqDz5Jt3n1uSIEeAn6wkz9vmaQcSbxLod0u3cWqbZ+/nT96cQIyI20TT0H/
fE2wFeIFvo3SDJtaZ2GKXNjMZVH05MTHCH+FuZbgggMlXw3EGAFATDDLs16gV0I4iH+edJs2Vh39
0dovmrcENO1KYRtHfWytM6LpSiQU/WUDjDX0P+b8FDQcWtF7Ve0AdwpfYsaJZa17ZRmtDqt2jagj
HqQoSNthmLSEpesS2degiynGBxm+tS4nrCLPxjsDWN9j+cpmb8RM5xRAABDCRIvC93pJBL5xJbjs
Znzmk9GcEadloJmOxsyomwybuFGDbvnbnKSG87lVVCPvlBtwio7uwQikNfNQyLZu4n0ug3xHaFAP
ejmKnzlOQyURZ2kIFpVod3t73AGucgqoSKsbYWz9SpQXUvaZd4fVdyeS2zMLDXm+gABnfl4nK4/l
VQxEXcl2Ae8fkTuARt59GJ5BcFGS3o56kqqrfETgskBm84y9iSphFKzwIGiYuOv/ZyN4dtoYTvp7
xEM87w7G2T085HHEIpSJWS939dHCLU+pQ9peDXJnGDxCqNguZPm537ag4zt7SYiX5lhDc9LNXPhq
T194B8JDUxiTMmcj7C46i4K324SAE7YIWCJqncsVePv1aCqvMJMOxjeJr83wqqvE9LwklUZ1p36E
exdtkKOKD0PipK+R6SsdqzqsMwFqjA/JGI3WKenF83cW8vBwUt5U5OCa+9bCy9pBNODjSy4lwiwl
Eub2EOITtK6T2gODXsGpCvPNO4GeSsnuNk+MO+I6p3MD748L9ThCcIy1/D6tPkqLrzTCO50cGULS
BN2mICQLuR+tUtCeeXNImpB4+66IrgoOx3H2Wm7se+vSzX5rnGbIJY5H7+Rew52MBsznZWW1Y9KT
1iSs7n2i2fcatSqaMnDaa5xMpaOVUptWaDS8kvkSsoXNjVbWETosZI61jHotf9+BQSfKKiXHgjji
zZm50qb8wYnlWp2zQpz/POJRV1mnvNT5dg2GI0FodNl6EMWnp8uLSzDwurtalNeLcXyipg9WhpG3
7EnowvM6vWtwuxNUzhuLFvMwBV4HAnxcGn86rsFW1CspKsr7jN2e8bG0AqmDhKf5GpHBa1Kcjwjl
oD689MuAOTPtn5FVy66I1y02j/K37HnT51u7p8WV2dbTeoQF3oqYJjhOJLpGu24fso0h27Gi75HF
qDYXsP2UYAEPx4KPor4bGvc9wypccWMyu+q/4x4WMqIz/oIzCbgVLDzFKOuIKwnZsVeCoWYu7BUK
zppmdQE4fZglwP9cb6BnAUK+ttmX5FEaoGY/kEkWsiKDkvYwX9kQe69R6NF3Mh+tejI/hnLTRXJz
tzzrLX32lRGnxnq/l3Sk7xALA5OImhziv77bAFk/DSc5lCepk7NUGBcdtyMibiLTptWqWrAkTtHo
onnyMymHy+fQwAFqm7R0xCbL+pXNp/yKy9LBSXp0ZLxxXrVDJACWBNVZlJm6c51qdfFUq0be+Kpz
S/kr2ImgPMCAlOQq40JakSZF6/V2iZRGDt7CZ1w1IysFWLnRxaD8juT6WVu5U6WBtO2s9ULClM+8
qbCsFIER+wh9usvz6qXwk8lNLm2bj6rYmksbtrFuGYH9P/VMUIRlP4bNfVlwBOLPFFJ+WE+PWV/q
IPmEmByBBc38Oc/XouDsX76qNLr3tLchgSfNWF8OrKtgSvP/vcqQHWfVgYyem8Cm7ZroEqXPJJzK
a1waO4IWMtcqq/S+LpEUIh2cphTClFUnMdK+tYqLkRXbTJxOrwq3ih8VH5cBPnf84atyo3Hje+co
m2sdryU8b3yrEPLwdlXFLlFpujeIlCv2bYzjVQK3NrT9KdlD1iPzWLFefTKCtLZnT2rjGgUoXchC
cy8P0m+/T5gxrleonsVDrNGXzgZ7koCu/GsfpzfNGeXKOrv6mz804REBM30PIWdKAU0YEYWa0r2N
fvcTH1GbcgCQtaoCPBL7H9ukPe1RYwSW5XVDQ5eSzVPZtGO+vFxPG2yYi57IcNI2tGZqz4A/5Xyh
GA79Kkp78oi3GfPW5wsYZs6ol51XVWOTHLRRF7pCaMUFMsncbYmxKZ+jM29Qhfc76TzPWd0gxjgH
Z9I4zbKjR87WdmpBugZvHhhSXIPldLps5QEr79177IYspzY/xfiJKkq8xrohEK8msq9ZdZd4z4cH
kVdqLP4d4dpwJqc4v/wPSNoF8cZkPbaap5JumloXXe4jIJIBfHmNd64TK0RpqJ7AuNtxjCaAtq/c
AQ57S97NhIGICmUzmLSxbZGMmHySLQy0citFWlwKMeLwjp704CHVrV+zfyQdmPmLcxqEgMJd1+i/
aSSkAsvx7ocsHBzgnm6rMWEXw2fggCSoI/S6hED8folycWyG2ZB26f1k5LQcL7Q5VwwHJMVbsXSi
kvhzQcP6MT4yjBuLsnx8t79LifX9hJAyUnj6uZ3kgX+dgmLgoFNbRnTi9ttg8R3atqsRSeBZas8f
xfMfC+hKCQyI20cQJ0dAvxlEjVEiEv4NwWiANpoUE+SkYFDdgcsXn0y8e3FMlK1YjKI1zwbjIaeZ
qke080qaItlsmW38UnquKprLcEY9hkzT/bj1c0I95lUXGJOTh7rtpJMm4NIbH7efkmNr3+9SMxqU
rO03pmOmnnsZ+AP/5AfhoRzE4Chz0ydtLXeppYaDO70oSjo2s8Q2kdAbv2dSP58na/VpUqN3Ax8W
nlfOUYXuEQ+9Ex81M5Sx8eaSTDP/d65bhTlJbYREk73J0v/8IHjnk+xFTT1T9LTfGU6KUaLJqTTS
sq7eNbo0aqfd1/BiqYWnuXxrvxfp/vPb7ru7RfBHicpVsGlx7ShMzntz723qn6acej9zJ9jMkmyW
9GKdg43no2MSWYQPvnvG05qJ8unXobzLsRJO48pYS126qxLeB5udsJyroGK+O5nGJonJeKCWR9eF
INFb9uLAAcIAxH3O2GHc7tlfM6kYFGf48lKvCcIx81k68AYuE4dnf+eHM4Fkt6SqYXEHBaGvfqB8
l3V6p/wymKLTyNJFsnCZSwkXNA6xZuEbEgmfuD+l6K/8NEFTsnrDFWKrEpPWX44CS0/c3gNEdKAZ
P4d2rlfONFex8mT+sZtooMb/ik0EqqXD3u49qqHfdghRjVSagcBYcoDOn4GqoH3K+7AY61i44bNH
GK4XRwZbRoTDh12EgIKo8HrjlcK2QquW/j0Q+0zfntkX+TrZcfhDUMrRzA5VtOgfY0tmN00ZrtqM
cIjVcx9SE07cL1gs0V8yECJUqVzP5YtQLil4OxDbyGWOen840xq5rNwF9B4PbCA7UiGmCLJFDeQ1
/yUSHVng3HWkcBZb8BZJU/TZjxDOTHx/InygjDhdWOwgWdBuH+SH3HzR1T3RoJDosWy0sksK+2dN
e+86+Sb5I13wLUX6B564uE0if2BFUIEmVJMTvtofHBdz6EsjL9STa/ZNfaLWbNkkAtF+XSvTfJiE
WdlCQmxzbSf6RjOH7qdwZL+B9jwbLUwRqDgLGlutNO/kGJv0o93UNThzpXPE4hJMiTOIwWwtGSK3
GtwYNjgi6+X+RJFgRVX6+6Lm5kmk7drdTdHiTPjYJ1yRZfxYOyAAtHYnIyqROfbpEpkVl1504r6s
/V/KLgczjehAack4osWkgfZNXw2jEXReWOc5MIcrBVGcNuwwYgXRvS5M6c2qno8a8xRP8ZBNDEQ4
xfty4N+VLFNCn1o0wFD+EZItEeXxl2sE8f3uXgnp6ItIWF3zYv2pJIcpJiFXnygfNB4zq+iyav6G
lgldbwrEmSpveIFCj1I0Zsvne1aFOP+CkE8H4uceas74oH6JeqHM+hVvewLd1tOthqp4/is2IEUP
0LZKcdOhmWEAjNzW2Z1Q7htyWUdLyZr72eVGp9A5yApnN199tjurOFgUAUZS59VeOgm+VaHGavws
BIkkWt++VGGGrqdd4PaV3S6TwXxB47S+ZJENiUTy0hjIvoLoNg/9Kc3HEW+81IBSjf8NCuubgyAH
AIulHxFaCYELiz5UnwJcRwmdgnshqxB41JixN0tmqxb+E4QsZHJ4/l8cyWnqgiOQS3EiDsIoiN0W
tSydHEf+pEgOtJk0KWXWw7/W7xvTqRIJntQdofMHvwugKqQEy4RiUlZqmoHSfVwRlBl/KzDl9fia
LXikx/I2a1wPtIDTbJOhR0w6pEeBYX2JomhRn5vXS2yrwtx6nLeHeSoTPOScYplQeWTpaL82D2fD
lj0LT3gt+fVzPm/EpQ3WoIwq5fTOHeApnUcRqOaPe0N/gCdFTbgMGH4dZMaaFHCHs6J/gWr21czs
Jme4NjRVdAfMQbSE/BA8vtTKJI5Njdz1/EipvJVPNXTI5OxCvHsxze9CiKNQ5t4EXpzruGIliQat
5aUhw82Kq68kelb/56EbkHzAOuZXVnn5jASQhWThMh4aJseHvORevIo6dW6Mf5NF17OiTCfFRPDB
44FO8SnMB14jZ3ZpnjYuS1DeTlIkzTzvvEqj84eXzXc3fS1rca2+U5w8XocorgcvLS8bHaJ+Ow3o
BdrM8qeePNdGA0/LItAo04Mt6vBhhCqKc4btsAxZppn48XKOcDTZKxj4/+cjOyPx1IcZiT2lyabW
NP4Y80FKBgYMlNP2GNMBFVjuioXj2N1oQlL3UEjSROcrecGrcgx3xn6Wi5Z1icKFPaurFsnMn1Vw
APmq8Z7N5FKYWopNcgb5ygd7e1iw0DjRBbGtgX1DTmYM/dEwezdnWvD1uDGTV5rScQGKtmDHnHEF
ydwKaNtOuE30LD/uTt63dvYdI6c7Kn8I+tZqqEoQYk4iEWx03StJvksdur1UQrznSzXzTNKHJlgN
OMqu3Q6X731Ioc0e+NseBQgMqlp7D8NnWanKedgmhQHD/BGWSWkSHG9sjRS98kkkCc5wJScApMxC
dQaPX0W1Drl5xmCD8rMJsyfqfG4QWnSL0DaYjDRkOkZUhoB+HqsV4xjS34I+u/0KlWu3QP8GK5qR
vLAFICayouR5Ycvy9CTXkJZnFPyWaZWd1CRqc8ta4+y2xyDffM9TdfUvlVktX9qanVVG4p6wKZd4
gs4sRNo9sjqr5abMZ4qWDo0t8eIeage6bEpNpVv2+N6U8ofytUt+FcqNtSlzyGjB4euVRXajItxc
ewGecsew4zFpBwy0nklPef4N06joVdMA5+3tM+O976ONN+iH4PB5HNSYOaDehkGzbBjywSBNQbA2
WIHeD7iAx9rPFuacgZyLWa+6xDtbETLGxn3aYYnDU/g1YtoVtdwCW7tN7Nq7NEW1oZClVgJq90Jf
Gi1OTKFiV6PWK6qQdIP/UbavMWR0EPG7MEQgt3UHGU/Vw71i7oc3ybzi6jE9EU4sCVJWSQuMjRSz
O+Q9nJ4/Wukk7zkdsCymcqD5q/uEC33L4VssxkY4aLHABC4AgrDzgepJalNi70FO4iwb6MeT6iqj
RN90M7K2uiOU7AI5c6XE1BMVB8xw27OAzyzFNWsNkpxUZT5ZwVYNAxQ4vUXv98BAlq+IYvYjrIou
m7qlaIrOIuPf8+qxjpj+HEwu+f7tfPDUYyN1nMmPJsJUJJNI6WwD0XZRDlKAMGeIFyBXdIZpQRrQ
YRcPUyN+ffiBmidhJN2AmjFh88wg4yyDSJ8ZLf/KY4Gue7d/Q5a3CBJLm+LXWjNUt4AYjXBzd+Uq
tMmN1lsN1MRhEHLpAsJD9/N61hvpH3P/W22Iz+LEF3g1YBCXSEUfm5yXLcJXtEYGV4nbTXamUOPx
WY5LKfLm3V2NMzVL9C5TQDCcCFMjKKWqpdJ52fwZ2Jnj52qLxLIHAvGBhCD2E4lVNFIXr63aOQKa
cZ3tITpt4KLicvWhCrhrSaiLoZ0Uj7ymsa/TfKl8xDNNPNGgltxW0KBXhAyICAXCIjEXIfppqlai
l2iWcYPSopaU6MFu5dyd7fDCpGn5koZ/wOsA1RGiFssUHv8AvovFJR5MvaVWxmkrPv+RwcC5EZLw
WNLKOu8oco2dfK2hABPruRSKA0yFSxLevERlXQyN1NyL0rX7zQHsxZteE7MHdjv6lC1tuSHyN/Qg
yl5lf2BioQdShlLKixn6fQeE3LJ+pOgLGF4N2qbLlMbwrkXiU5sm/zeFxuEMMWM8/SY52TySSgFw
q0LaeaZxRN4iI+wvIeMWaJtX/MSnhhHTkh/88HZMb/G9VGgSkQU9zDgP+FEsz/Q9U4j0DZ0TxsAW
OKr56cYsDwSpiQoO5OTZdhMys9y7BIBzszzWlunJ8lO9YJKIChTlTuYOQWWpn1GtcKR16Qhvdshv
vgnLV4zOJi4AlAI7fzpOVyjiZrZSHP2gOxbKy/4jc+S8EVNCUSeoD+ijVrvLMnmB22JuIV/sNKix
/1/aHXPcgZUEvthw23HcFUBIfQpmgtACsQ+EH98wORxWGqZkOmi6JYX43WE2BZt9E2WFqKGq3D3c
Suy2UHT0o2Fa67GZI9BgqP1Habq1GaVg8/yGHHFsqVODkCaVbw8gDtt/YdvGmojCEhGrusLrzge9
6/tqNZMcWL4xZtkpQ/mJthgBF13jlM4OjbDhrI7OHYSOTjoDm39Yx90hQOKt66nVJ5sEVSgbpAvF
pP02B0P008PxrZ6ORM/8RrYr4h77QgVzaFjM/safgStX7gXbfuF5EvM6fwh7n0seyCgkrHBqNvZl
AO0hXg6B+2/Mrriam8eQ8dAQJ6BAoglU7Zomsd8gFYKRj1HINJkEs1wQHMaJcdGrTzVs/FInOi9l
SUZdUeyDkDwQMv6kEHTIxc04bWmw9WCmwTP5I3+39B5UBz3TpCn5tUijX1M0R8vLDDQ4D2wu7jAb
fUsaa7mHDMkzPrGIuO3ifQV8CqBGElghM4+XYnCOcnCQEv46UeuLov8PAcK+FZ8nPcVS86A1Pjgp
UJ2Bs8+OSprAcPeVQzVugFf2EQ97qXGGB+Qv7CNs8GPM2lAMtjasR6Ann4Ag5WgFUiGaJGRz/9nQ
1a6duKIO4V6xeA2sSRFC+gxWOL6MJKhex8w4BjbJIoDElZtd1PY6wzN6KfcxpmQIyRQ2UvuL/Ck2
1MPoWORHsE2XoCa7sRseDZZ0TilDyFypFcnXgDguU27dminQYM5L3AAUDH4mGN4OIQph0SvkYkxE
us+26YrxfQ++6MdLBl68KKGirMdVTUkMADqaFtAAlLP2ed0vXCNewMkPyZtgqC5R6Pl136NlXmn4
ZYdVqLgoFFLgGrzAR4n87yRy7OS5eGdSNLCGl+8Y7Zyw8isULNPdM9ufmBLLg1tFvRpATROGKfFj
/7fHCBcRImT19w6RdQC+8sISPixQzEYLF2HP7L600JV4nYs6xDwK0FRNABE8PgoJd0OpNBYmEvwO
ofnJKV0w8eN28b6lElHkkMwsLPzdQPhuLRph+TlPdhAKkWnihcfOlNuLEVcEtrL1k4BuUiFMf5MX
yy48FsDlrroioiLWrnARoBw+62pzNKeAyoyeSt9wH/u1LUZYlxifKdvuIbh+TFO/3T7p5jNVadVS
Fj4OPIUqRT3Sjn4BFQ/tw4baUX746KdewyoNeEBVErYT7No9TT3B+7TDdPGmCeBSniprtOOsXsR1
sszGlSFsrQkblWpd9bEbY5bMHhMNaISptk+DV0O6/k29RlxQv/XTLxFqToL3CBGWKv45JMd8H8bG
PXn+Y0qohHpAEcBE31r6OwJl5339x5AHV64O9877sF6784uIrbein2mxClu4rTi3yf1dpjZ0yBKR
6uqood5dvurcF6yiO3yXlNuVvd2CLKQ8lmX+vrD5iR+hoQIS63OMJCxdt47qzswKBwM5+EqfSd6F
5tAnxHFVNapmrYJ44KGADsdLthwirbxYH74NSo/BcCN3qMRoJLlSepAa8lVxx0NN7xqlAUx+4U0X
jTp72wfhvTEApN1SF/hIUSA6toqKFyJstlryxo/jK4/zfremfPi2OyWUydh9uuMqYF7fF5hkL6fr
r+9kPBMcm73g5AZ+FT4DGmlee0MdMjhdoNqgtacs69yMd00sFMz7Ua/AJYucvXj0Jh6R3i/qZBNe
RoZAG2sRxOHVW2JrNVpTavf3HJ9PBGpmZyBLRXB291ILpuTINHVymmaeaK4lDaP2nvdgy6omYuPl
LPfTWLDpnv3dXVBN1wv+PI7sqDfxtouXjEEkPBpuF8V5Namr8saKvPDCc/MXpBAqBl8gaON0CiJG
Uw3tnCC11mwVynlLWo4mDOVjt5y+7jSylVuQljGo8mPJrtUJKSX9xNy/b20yT1sa5hE8Rnzfq1iM
3nj1Y8o8bIqNsfalveamYT7IBPj+XmGqm8QQIcJeJRRN3VTGOSvBD99yG7Sp7cJ3O8Dmb39PrhOo
YNttA84BJ7ROBFN+OWKNUZRzxu3AasFXN+XAXLT/c9/Tj6Mmi0t5R6kYshNFGHvlvQhel5c1v5U3
lNS8rPLYxZ8Q/tOYJOF5SHydoNEzUh1+4D2xPAE9EqHjsvH5uyDbB4HdjY3e9+DfAk/IEcmQdLPu
emtlpHWzG7VR2+At1ktj9Kq6keO/bsxh+mcpHjlyVDCQU32YPYTb4qeFEeuww8bjVEZcT5INAk2U
Iqvyo+dmbhYb8WPBcTPakhPH/eeEbw+B+ugLgn4pdVUuEorT59GjqWa8Bg5Fu66SaPha++9BJFlZ
ZJnZ8TASUvjRChif09OIlxEukzNUZFCUHBON9mBk2+SAM+szfGsZ0E/n4/6C+jTHsefzrTVMM6eA
U2Yf+KQB03w5ul0EUfNqV1UTaNdNTNFMBgowfDnbMEFwh5DXTZT0tbsRtOIxgF1xQjbfukWKNUj4
nUZjVdkNJbiRTbsFJUzGKRhmSTbSy70jcZiqhXX8jzx++v3ZpME3a4saGWfkdjQNjJBJiatplY5M
oi7QxM26ksTPsODLHoBqq15AoybBLM3s1z5cVYLSA3DgmRJw/44bEM/dvnFiKYU1EwVlSFkjxjdH
rvdLi7T81VyotGbHICz3Cr6aARHEAkT0MvxSIX6JzVIToPcHh6CIwoCM2TY3+xi7bKyNrZtErI+0
7i89hl/p930UvJu2o0BTF+P/ERq1kt0hERluJwyNKKxo96JyawPIGf1YCYnmyBJiNNSBfslzB+uE
yWjxRXXiUpdn/khAiNT9+bEFEZxpoLmiLLW3XSDaaNik7SoXpRVU8C89y0kQHbtv0BJWwOmY9TZI
1B1sOqkScZDtjEDwVRBbG2e34Q5Q6DDGBJYUVsBhiFvy6Sw9J1QqJfot8ramcyUHU/09KH/gmIgG
4uPYjeDGHNfSnZga/g0pggapIRqO3DkhJhNIxRlxYmvnZMkvYZMyYXxmyo39ATt8my8gUnYLpfNx
jP0Qx+ymrYSL+/5sXF7AJMmb4byaXtCwmVHj/8zGPSUenhK84YuvIyX16yDZVqycH7DIalDfJAiF
43nOfPlYDrinaY4OKb6m+Ea5/PjkARjfywxCNTYfKsf/JFEJyamfhTA6o9y/U//1PDOmoNXx5rz7
9eHm23iEpmzMRbOyC+c1OuZ0G6o92bLk7+TZ2tKZQS+yQM515gFLrkQDQQjCMaGsOd9OUggqrDiP
dFo5He8zymwnpINL1kLm8Hdc+PuoHjJugKl1YvKsLuxrTYkmW3B4xSjuj4He42tIHTqNNPSBlv71
5TPbf1Jc9NcJZyKtsYSJiioKvK5q9DViMC0XXeWyOoh1Z23TfeqINUZLWV1l6b7B1A2s9gJG7O/3
Wr0g2soiRF7tPIPUyyOike6iEmpXyhZ5B6/n3o7x5eSF7PAyCO2uCWakPwNrJFEG2dz71BcsK4e7
tFVrGsJr7PtazV4qyQ3kVVoGarBHUywByG6ENcTEeAShAlGNX1ziTl3Jt5hnBSRhW9NdBEbOwBh8
ytgE97agXx0Ympy5OXU5CX3PmMXyhZQwMZIDAP0YYpLytnZ8yTJtPJUVBoEWdf/b8UuFfQYUThwl
n0aZcdOjRH8BogaAr9KoR1/6h3pCkxEaTOhj2nPmrlzUOOVq8YDt/4fz6UY2TlBwutP/O3AATHRP
RRVeVasm7cllALYO1NZVAGDkSxn4zSxNLRPB+bzdTZvVoFJB2e7j3eVhPIQdVZshFgbA+/Bw/Aq3
aaTdFfG5XtGcIeFjrKWHb7HtiWzTxlDQhrMsXvulqGTryp5rvvJNfrrd5OHlsEisyhvWr2S6xW8d
zlaogdNXkDpKXVbXVFzvnjK5kSsfZ1h0BnYyh9VNKYfHs2S1g00BmmYR2VabLyxbCVLjHKxG7+6X
fqY2Lym74A61v4b0uJYzxu9lgffBII5ERvMNNHzGMc615+7sCeaxOGDPWmAuwNTRkno4rroDu0R4
0nLbwS32glLZBykFTuUwvKv7ObMu9v38JGqsmjKwccPgxrqMlvI4yZffEPbmkk6O6vboI2am2pjc
b2/PGIAiIq0CjxbgiCUDdlNr70Hv1o2HbzMCJotAvPHYaQNKuH9/WfWyJrG4+c5gU7i/QA8cbPJG
eiKV6jSCqzybyfKC8DuGZpg0wy/2Jjej3Ykg/djusfxZQa6ti1KYdxQYdnSrcCB0gmnYHwRB0ORm
Czoln/qGQt5cPBFZCe3n7ScmKD/1Wcs0Vn/HX6HNWYJuxzWsa2ZDvs0JR4M/rGq+9l33jG5OPMZ9
L2mlrxCewY8Ven3TJlp6Nh1mFiFy96//Fnn/j0Yl8gIzi3wZ+4OxQQWx59nLs2u8Wu50D66GV/1N
uIX+jI7ud0XKWOJNhBop44EAUONf0r1LnWurueK3WcaVntOeRwow92zNIRB2RgdzdtzLfrruuHaS
6d15qcd3wFybKqAF0MREf2XK1gZIAuymB1tT4g5krWEq1wol4Gvo5kUjDrVJbF0CdTiQruma4M7L
aY/OCPMiJTQWZGl6ZVB4YSI0PZuOvCyo8TRyMXApZxL8c9fJduN/eX9kbjOztHaUWtvFB2knNIeg
QCS0zwS9lT19UtJEcKVYdQZMB4LCYKymaCyvNCD5Qk8Fca2P5iPA1zusd5ntOYDihi+ye6UBHEUS
abDr92iqE8cxgx0hiJLl19SVP5svqR51IHuIh3sxpLzQwBRRpI1HdVctit7SfDTXJuv2BRCkmOzQ
Zi0qAguM2VAoULqX06AKiB/3Nz0FhWm4tru6G9JMdjl6YBqJhnf6gGzYL7K9hFMCSYmoeqMkK/F2
4VR2LIDyPtiF3Gh4eRn312PHYcWy2NKyVmAEa5JFPzTEtlqv0eSy5hXtMJJAbcEgum9DpaUSQLIs
41bJd+lo1XnY+6Rdz3w96Ul0bgHyfMBdmF3LZdFXsQ0D6QUpOUPEtMBOep4LsBvKZrFMhkpTJeQM
d6KxxXjIunsQhpyKqeR5BbN2x7XwbsxJfqH67w1Ly/6LrM9laCA9Oi2ZDwJ2f+edpV/wZ6bZ226f
41MGS86tW6RW5WU6Uh8C32lqNRhHyjW340Xi3jupmnpCMgqSc9VqxeC7mJyh8tnP3HoZlt8ddJ3+
s+x2XkDkzeEP//NZEdi5xHhTMWGab1PICinzknfS/o+JAyjwVd//tsZ9cqbwERiw4fhmcC/76vdT
rvlc0ZDS0UTk4iHLVYGCdhq85lk5Y6PaGEKW16+0b5V/GeV8Iq+5Vx1XAJBUKp4htc1Ur4sXpSPM
F1Uo7kDanvJRaqNr/CO4MlOImGFJmS+MJDBhVLKWkKYofwOTAqcv85nXUnX1EA2Kdacz4KhrK0gg
xURO+QH5fRAjZ3sP2Fi3NezxYPRTB3XFLBseP78ufq0EOcFD4USe6RJRsI8/G9HvGrb6ktwATobY
HxfJyQk96MlRXBj1fu4lucPTGn2bewV1nzbLbwQwMiMbnpkuJsTIMFC5vfFtDpwfuMisSoMUV59S
7HWNfQ6g+fDykTd7rdBCxZYhC9Amu+nCd5NWj4Vq2QVUgQKuBxW8oOKK8NICBKH459zbdl1vmCzi
LabAkOrf333iWggkZAGw6J6Cb3vWN+MNMt9La+zABkSA4Ygx/YcKdzrBoEcMfSm4kvTKE2z8DVAm
XoVMdVbH7tkNCojLip/3S3RRzDt21XVdYZQF78YHexyyrPUGeU/S8LMGXMDTdQC+LWAo2ya52XpC
pWNdxSEarSQ+97fGbxlm/ozK8KJYCV/6Gegs1dDucpW5u2eFf/97Qbm0/RiiMjOo0xGjIes6eDY3
Enx/x5yS2S9Ru78KnGSxI6exMfhKHbqGPFgAQP4cOxLWNFLRBjuc2DSWe3RmP5aJjqxCISJU5aHg
UM98QC3ZMQ1gfyyxemcePyPDcFHkFaTQOeCu9Hnx1QCLYmD6wh6yRMP+l8yllqJHGBdtz6r+2RcX
ChNoXQ4S/KDy2rPghNu+2ELRuXvljy8rmoVT40PdqokNZwEOqOENoqFRcrWGSqgbeVs+8PuLjee3
9xQB0YJD4Jh6CPYENvjxCIVHwbjr8igsnU7y8RemVwalSQqTXeVCIJEABGkqXh/YAM4eNNIa9ALA
Ldcn9LdvWlEKcGNfZ76SG9ZkjK/HSmp9HgQzl5573X3yGN0o9wGUsTF0fZxiwAV19gNpTQlLsVM8
Nx4j0cx9nMTljlCOYd6jlivMgPpxtL/oVc7o0YpY9gTJih2kahc1th5acnSS7aml1DZYCa+4HLW4
e6e/ScIcK9t4tA+DMHxF8Tp1uQzllrhX4gOTn+rAqov6+WyFXVCOeAH1hRZhimVdhoJkMTNhnWFM
7CAeF33JFSz8KiVtLr0Z8h6sy2SXPdDCnvBzbBxzXbd9IFoK6Rk4hglsBGkTRRICgt+6F8g6jnZP
gR3nDWnMH+VuAE2IFQaIrro6ViR20OIT4mcfR8BZdlzSANYIvFHJm2PVIuj5UPCe+FX8uh1DBK0V
/OtfxSZrChxxLD23VpljZya2R44ZS/wIGKeOQBGS0WX61//b/JOwQ4iynG4ULQR6X/dd9oX7fWgO
P6Ta8FqIrEkNqryMMo7UqpKkmySpATj84yWnFaGcg9Phd0idOG9LVtPdl7uW05EWI4QOMOpQ4p0i
SvtvnGc9nWtoIEKQpMLeCjFE23a6QCcMHQuGOdFCDk4koiTzdhrCagCQkJ0StVA/2fJ4T9K3ji6J
ryPOjmJyZoy8ap0lRIs/0wref3H5JHZnI+2y+IQc6vWsfg08Sr6ZBezgoHoTeUQj4Vo7eNWonF01
0rcBM7NDsmVAO/FHIBvuBN+qHLGUZknWt45vjbziyDV4xyg88w/tslYJt6CoO/0WTWwVAVB10zO0
GSPwW/HEfhkNF4J2nawNC9ogbnsixvSqFgJ6fW0CJqVwHuhzCJerBSYwgPFdlU+93CdewFEqdryQ
Sijo2fXgw67f8ZnVgHj2KJmKn/VQmFIgNG/kzdVj9Uuu4ic194L4APwiCarJWyNJ5gmoaAXrzBFZ
ZZCZdCqev0bQIQ1xOhz1CMozbHs0YNKZhE8ubehcqycDGJikhlYAqJG2/CVQtUvW9tiTwKxD3MfU
dSKK+UoaU3M+wkkVuoEHb75kFk6y56NiXxIXeAgJy8fm2FS07fGTzXCAcP7AReMNYQaF+NN+SHMs
1Z1ExUJ2siZp1MjsYZ7ID3LSdghJSsKTAg64A3AWhZtAeD8q7+kxKlarn6Xo8pvRrtWMP38uP7Yg
qVKi3WWvkUvnBWuFUe+4JVcPPN1RBhihXqK9sNvufMrzSNJqr31ER9r63lBuxDBikAEsbNoxFlTy
gWtylgAA87SENjn39tBTjPDk/8UIl1sd3uyVj+6l9+au6F7jes1mgpka0MXVVsfGi86jxLyN5CRP
XMZuwjUmlqfjkMAzh7qoE6yymo/qNXEtIeOvfYTRTgdoTHPoCTg7+M8OFRKMPP2GPWyyZRjDCZ3q
GZtI8DuUoqYCm255hSczKFM6U/CjEHTDBNywE40YPJd7mDSxfZySiW0Jtt3KffUo6RHWMW4K4sh5
U/62HINadWGGSVezFv7U0fuGo9I5PdgSw0oK3V/df3Y5IqjnIo4PQ4ET+SzNAKkjMxg2ql4iwKlC
IZ0yXgHhi0ZL+FJEKDZKZx0bj76MyK4aKqr4SkpPL4fVuhW2Yn/zgrrOYSJpuknNUEoyNBZ90pGo
2FnikGTRcEzi9PACt5OJRPZCpmrg1UBUk0mvcGDJ0SdYSre3Y7LVfDggk8xGojfvIvhok1OfBMDs
vHja0Nzl7ynJUEkhwJst920fQBAPEiDL8LbbOWJef+MjStHpXShduasLSAj9FVMkGuAuYLWlNnDS
r93P8T0kot7zhy7LL36LUKRNCw6K9HElEo9VasR02XyMAql0Cy+fbJ0pS2Q7x+r1KFW5cviGmhDQ
Tdv52gQfq1d4VXQqnO2MgapiOMIJFqJygzMyFMEO2SdkdT6/CHZGkxUaG7CM/sN3QgkvU0eraugg
ZGtdsfVhh/qWUIARPuek3pDrz2mLtW3dqo78T421Xr7YfsmaerqGpSEoMVjyKrhMJKuX0FsvAEWQ
uENvTbcnVt7PH10OB2C3pwN9oyG6Y9s6nh61r74cj2wcx9/5IVJcSVY+CXX5ScuKaLL5JC73tJAT
D4c2+cIeCjMpXqvF+qqD9Q4wWzyNX7WwN3GKlHihBaVFxm3ndDyCBu+rtHnzvrB2JfEQAjKsPMpI
ptenw2cLxNn2fss8ZJCv0RWAkXX7NLGnDtv2QDzOd6CcGUy65wb3Bo/BgmjLoP9XYWzJCwOS5B3B
Jit+tSk6b9kTSy1Gg/DrHzPhQOcLuWTqVhzH/Jk6rzRek+xP0KXUnI6Zt7BhcN4ueUpyfVeWFRvj
4YvVe7xAUFLosG3l5f3vP3Q4h2zkPARCzCSekWBCHjzWWYQFFKbKu4DBmZKujH++4AMp4RA9Ts7c
RWlmg/xyiEf25wGcR9C3jNEKlWbBRsGcLPOnLv04rGoW6eMWo1yauQyJAfHsM/VLEn94/r2RL9Ng
d0xXXmTq32EG8aNDLSAf671/0YvI+5OeZMD+Fip21Fd5Sv2b19f2GAgHI5GAORGdHFTOy7EJtQlT
xFuxeAu2UyHJQVcYSqc/0AyJdxSDQBqj9cagwjV6Muofp9+odRTsczPHMoW547/zrG0Njlylux8T
u8OLomQcymAX/ZCBUeIID64OcgLryEKHXjkPZikgG91AJQroGqc2cOISCQIEK8ONdIN3V6ADXKG+
PdyGjnXT61a4VUte0TPykGzlad6ScR9WqIHhl4CSvHfaGVIX12iLyn5ytD9luZAp1lk9Jt2lrBlS
Ugt0vKQhEgbWadowuJx3RzVo+7DwB3ZuB+d4IMLDZc92N9N7rNNeHr9cc4wRvht7tmwXR4Nt4Uex
yhg4Jp0+d8QzI4rTY0ANqJmRaukpguBPc9tzs36isH/q/aM2E6z2Yx73vspW8W76PEJrAhpRqyQo
fjAtHH2B3GS6ZQd4vo9D7lbl3qqATI+orC+J5BirmnMEtWvcwThMEkwbsMeAIZx+CoUaUFODFFUg
0ylp/dY8SaLw/r4tITcK353gwckOcnG/Ztc2zAfVcxdrvBSf8C4A+SWg1dAZbuQPgxRncIIuUrgD
42Pg242qJg3xD5Z+Task+BSkz0OMmp7OJQ3vBJzbWSY7Xo5Gg2c5wtWpdJH+0+XVaPsFwtlNdPWP
HTkIuO/kkjO9tM8q7giaFbhc+55jBzoN65oDUuxuGgHFNWT8NJQ00lpQZA3gdmSR4RiBWdIlEZ5l
ERg3BUaE8bsUPll1rY/EEfrlkZLngZNx35ImTdfoAOrm4nWCOc1ODj08h8T+rFGKZWbT/5xu/IJX
jKcOJrWIz6OJxZnQokjTXI/3dbNydUNIU+fbY3Gzoikfo7Br/pYxCV+pHElkG9HllAz1sVWj3skR
mfSKxL8dmbWQ2LCpE/Vf/ZOj4bIzSm7F8ZLGLQuJkS6xkqe5JMdyB8cdMKT40OYZ/znzwHRMZ6uD
lLhjdsn/ydTK5wwPFKoshaShLw7YjeSD6QtUOLY76TEP05GoDyJhTo4ncYul9ht0A25+tSTH8gcE
CDLxmGbZL9vGhKtQue+ozDKJWdUkiXRvp6bTkBIwxpn5Qe7JlLX9tkhSvVSN60SuM9fMFZAfoF1R
8IVgGJUcdFe/34yW0Ib2i6I4X6I2WXCMNHJUac4Ax8ZVsuVZn7+ltaLYAO5P2p+PcLV7MHiWykLV
0KttQT9uVq99/ibwZJwJePXNoKQKL04pPmuSA8M49Ua0oxcclkatZuTEQaoTe8uWQuhPWGLAI3Mv
1sH3wh0uw5LUsW/vZxJi4jDSu+Dc4VjX1u+bhmEpapnRFf75lADuyheFprYx5rfOeJUMZExa9ib6
JFwC/zM6zYpzssO708iwjQfwgMErUgGVYyAbY8ESz7avnM72ZCdh1eUiybtp9lRgbgXDfVEzjzXp
zHxGLH+cLsFg/FJqir74KaDWHTuZXiJmtYF0snx60o5VEMvRNYlMfoK2A05XE6OBJXpkf44SUP6h
y7C2RNqHe66DbkiDHVZwQ83fCyhrwmOHeCxOz+CA0JqmUIymsT6X58otF4Gl+sngE8VEYDOxrYH8
UE3Me489oOugNx0SU0j7wNIxkdFtk+RGU/EwKGryYwfko75ENNpHtfzD0lneazE/fU+5ufv5kks6
F5WyX018+QDDke2CELwuVhM4AAJQ8DKl+DYYrkv3HiCNJjwJ1gHcTBdUwoG3JfUruN2xgIkEF6dB
ApZmp7Szf7Vey7BqFxgy442lTW8X7kG23NOMwwnqrRlal+S2IOg+h797Mbn3PxbfWVZkbuBNOpJq
+QZGRbjeLa5Fl1Mz7/U7AOQt7zBF6i10jKt0UzXuX9woUPxFLAZsB9kTNTv8vv2wk2uzr2Dm9H4Y
rnwpe1HxuhUZLPt2Okp9pJ4H44+M+WAIG3bBJWE5bPaP3GOHAnsuIFV8ohPxMuG7RD1Ka6V9arxf
q9JY/XPyVOFMlaMICYENwS9X0evhScA7CjniddMi4z55C2LoXQmjdbMQ5tKHb+ucsOJ2frg90/Dn
MNpGS/rDI8CcUqjdoJR4Wj8CEoe0VeBLpwjy+ISSW/8sJ2csY3AWQ5qZFUSFepPTAtycUe5NprdK
W+IMVpf4hu77t+xmVBG3zpdQo31xYWvdDtMJ0KtkddLdg7RaXk/JX35LrufQqbOC7AysG1lnKDtL
7ugu6Mm4kaViJk+N56Uwkw9OP4ToTRm59wyTg+Lx+7Alxs1N+Rd9zRRP8sQHSMS/S9eg5rs878rd
mWadaRaCTkLpGxwGVS6JraNn+HLv6AROQ3d1nOVzTWJnSgfBihwZXcW3h2zF61d80FZM0GLk1AGe
bdcoUyoAK498l7mE2EW1mvBHZIz7GZSDfK3J3Gjqp8fG3xo+oTgipfmNqG1sV83hnT/XSwz76oHe
dJX9ekHUMSgdZ9RRscKg4Z4gYWiNl0Ph5gRtQFypNP8qzUsNIyQXpIwhYRSrvht+LW/6fqK1UpU7
djF7ftYzahJbM1yhyZWypeJm2fhp4Nl2TCb65v69rbWAG744S1uvhEa0YdQlDaOGS0Nyzw9zD06/
+gsj3B26RQPE/6cnlxvTr++SRDQGNADVLIuC+YUuxHARBoRo609r8EZjbdRI1KBcCFDbBXUZnDBW
A3Mo/gCO4luC+6x+gyJoYMp3y+ZOoI82yISF8H8+3TUiHnd51wktCmGDrhv2uyTJ/659Lcjt3aFG
3NWt+99PMB71/tngCPw2x8UC+/jUwwSR+8BJfgSpt7xh5V9VbtR91fqzm59Emw+GzVnOfJyolTdd
Q/j0UsJDnbz4iISb+3oG8ypnQQXi2RGjkW8vtAs4XGzpOyjK4gNVR6BUhYlBGlmmc6t+lswsMrsF
BJMQy4Y8wMmEuMBmnWpkzS+1Hk+agVvu5F4BFtfy/xMCoWCHQZwcPXb71jHGuhI+xJRKu04tEh5W
6r5O+/GY4rzFmmwzVL1DPMJwNdip2r3+dJQaIGMcjl434K4P/ZyqQgbPYiYKq6kMhdGRQ/KsT2R9
ZF21zRLFdHNqYkRP6DKWAF3PSv+6jE/WlVrae+Q3bZ8NIn/WvJQpjPejJRE5hEiFGobEPeeM4sMm
IWCYBfAOmLYKR4RCS1P15xGuto97rVkgIUlNZvnd2VrABlLcl9p9Gw1TmTq7rmGEnAUmZH7Dg2GB
7rMwMOTTZL1cyPPsP9O4jakaorAqk9XDTYtcTT1AXknaKi4bHS+oRFISkoBOXVEbk17BskNhGur6
QrXwz1JwmnRtPj8iy1fUlLw6vb8HFe3u67gn3mz4bZL7oaIfIL/FxoCPVXsvioqBViXphrMG+qRi
LM0QENy66XMBMfEH6gFJCCjV77447QJaE8nCSdm6gPoEp9oOwHExQaQMsIFzd4hMCnmKF0IDqlgW
CBH12yToSsS9u6aq9lqXK1k/anuWogpSxPcIdK8IbBb/oQjQb7/c6+WSRT3Wvvbey7zKFWLv0bW/
S3f7y0Y4OilTGLXv8/WhhjSUJgn60ULeN+KRP386kwSiz63hJniXcW2R+IloCsHPKuNTOysFSVof
8KuxILnv8wa112ziykfcHe6G39460WH+IIUN1E1QKTjP7GohxyaoAAOPjca8nzCc34+gRyARciBV
YcVnpXrS6eykrKIrdAnwe9Gx47EfOtb1gZtq/fX8t6sYGfLRcnh7SdZJLt/3LqVutUTDkL/OHwcj
2dIff96jn9uTLecGd+CuVCXTP8keHcjyVHx2kI8EkfJsXbTFTWX0OsUWRErUAOiwFcGntYKst3Oc
tOpDQiC2S39lb45KSGXKp73Y1oeDXBTiaIIWvU8Sx1QGAokyBv25MapeP1bkBN+zw4o0QWU+fNMN
/FMuCu0gpVBfU1+lG7M8xiaxER8MXE1HGZR8Xr6KK54X/bqtb7EQkgUbcOszLq7KE0gTJhJxz8Nb
aUXQE1yKQqCMhtjOHaffRCqDZQXZH8LngtJLDxXWxCVfR09cKoiqCz/2k9Yk7kaUOXrscp5ia0JC
hjbisv048YaBbow4lEYzOfn0q5nBZRTY7DOdVR82dptYdO49i7sBKBaK6W9/xsVIDxSFLAkcTQ0K
Hgvr2V4qbWUfFEjvZwXbCSYysMrM1Wjyoi5R6a2q2kqw2JnyhFOuIOPgN9WOX7O0aLqDRXCHBPGp
sVpOi20UQdo4DgGuXhpDDVjXaOpNbyQPqI4RDcXO29WlR4IpeTq25l7RJ/259c5tNn8XG+0JVNiy
ZDGbac4wseMQdrxhavb/4Qy4250L7Yeh6wTOwYfSOMeycq3hSGbYgc3VUZ2Oht4zkL0kigtCeF5x
Vc/Cqn7vQi3CnbTgGyPBXC+1crRO0jpmprhZr8QNSO3Yd9f82XD44tuKJ3L5n4pNSVU5fVs8Bx7E
m9ozPF3ls+FbNGVuYFUzi+zLtE8bxIPHZiKn/xFuRBuyrlLuuaezq4YUZuHuSMDnZJqRuk+obi70
y+5D8uiuIv2BT9bprKQOWAlxugDopNkHqIIuGVtGJJ1yTc0+x2mbibLG260XK2kHyHjoZiZFuf/m
uKJ72WelpXM4jsOiXraYrk90P+va/DrYbxZlERyN0WxEwXgp7VhIf5RgSelNBhCMoVA9IkWCB2Qb
wHOg4he0Tu5evsM/UuH9+BSiWz9FQtdcoJF04ifEbCD1aLgl1U5VA5J3ASfsKOBjd7WTe2lqeQ4o
8wuIn66XnFCDg/Nr5aSsZ8dsMu2/yTyNYViJT+nBrAWmYaVJssxDoTjNOnZep4wfjV/B6nh5QvaR
LndKVcOhuIuJATl1ATw3PAtNmSv+HHXmc+yaEQLpJWUh54v0aKWFtM4zHZ1E8C+2XUvQ1tVHPOAd
2EiWuTtppQzgtCGEp1OHFg1oVexqBU6pcN9NqyLeDDNuM0HxyZd/Gy9bvUoX2D2NZmm9I+yHsOmd
DZ+y5sdhJnsDoJPPxtp4oHwB6LCH20Il4OUTWHJxGA8sPBiRRVVmXCwZhFeWLxH1+wNXGkcUwjHl
mOSqk5FPJdhZrZg6g6E4yVFsjo/FdSruukY0mytjhlMGAY7t/g1gqYme++3ltmknbnsLx+J9Yakf
jFiRyy98+JLlomQM9/iZ05F6zUAnzGIHn07GdVHpigxM+XABNQrIqG6Q9W9oJbKjQrLredmNayhe
2ca0RBLlGkWh3lb1uKC9UAg7Ivg+lWMWjqpv0gtUN5+t/Rcg9w/y1y6GMo6tjtdb4+ZUxwhRM5sI
SxWBEPEDNqdD/reo9a5m/ES2My4fT5gZ1gMmEnl21UPFtm8eqMIJoe0KtR/Onuq0oDbJU0U5qvFd
z2GArIzlDCRwZJG/4jt/H5FzLnIV2gXLH+qARhb+htMAUminFO5qGgykjMJwBfp5KFPwvb8LHlmj
StpfLJukuLko2oWWCvlhtBU4h+slyjEnnxitbmp22JkvnmYU6RXKWnn1OfrgpsH+zFxA+l+wHG7G
75sJLtFjR1S5yJzSMpL2G1He1aIcpvpG9ZJ2b31A+3H77mDkErMtSBTgVkUxbt7mFvBkRk3RF81Q
jmjYgJ/iAGtEeTb/67gjhtYx5sdhfeWYZT3WCP64vcykkjEM/Z2rOSAJ2FgZp9nfReYvvdGImKri
mOfwF80JVh8B1RfH0kZ6eTw8x8aKyFK53PUOOTRzBCu8J/+2ONvSW5GrlB8r83BTGQZfCG+FOT+D
888RomFNydFjRhWvVFcJAd29AJScePTYFNE/rxWvln3AVU+H3fw7YX+i0Nz+/CpuMSAcW7jUGQY9
6nsdFO2WvKCMTUL6vJyDujOl337e5wKDUPfMarY2GWbxdm3iYM5LkIW4L75i5VMGhpGHnUv+Zjcp
NfRHdRJ5WszeR0WIDC9kKW/nWW18qnq/eF/RTtbkRoRG45WMdTgVMQVFhXQPdkXiCU8bOzZaZZ/T
w9QwCfoIO/4RqBVYK/h+akGhxnnoKkBgCRMRCq2PvokXS7dn+mbhuIErOhTVLnEONexrb/rfAEDY
r4X/36GoERNA1ecVcoQxueixPkFTcO4lNshunQng53HhdKydSGxnSgV6wIa5LyaLkESP30IBg4pP
hWN5wue6yqZT5BZHIoQopiL+kLjAV9XprH+0EPSAypXr++4x2b4N+XaaEaUZkCSeD4wdDjQLqBc5
jlwA5cLXQ39o0IChets6wC6yqp/8ow0wqstDrZT1oo+qgNzL9gu8wwJYgPKaCRb8ohYkS3n3oYMH
xgTPkT9Lr2U/6uQ9duHXsOkTP98+OwHxzO1lhnhVL2a0uXOe5lN+YCFCnZN/Sld+kWI77oUaG/yA
zAzvTJqrTXO024uP57osJzl/yQwdCFuUx96JYXb1PdhHefQVNjjRiI4SIEbIq1kaT4XJ9Jl+S9/7
ePtTDtOfqeexW/e1W4Oxtnywvf/6GSiUcjqfudqtNkZ/LWvrFJ8sPM+feuxjcXKDGRi3o8TxPZLO
ZLCIELJT6Qy1MMblOEVb/emwU7OIsS+lTtO8LN8vYqYQsm3CrkAw3XP0QHQKWmxkaRE3xTw3f9Qf
0Tj9hmNwFX/EsefCMu01VY/KDnoLuv8lt28hlZ49VD9xJ9sPr+H/0E44HUnWVZnR4zYlrUm6ll34
wnI2TWsZdaGTJZzW6dLfh7HlNccXtQBa+iKHJvYIcEgeRqtLcCgL7g2kqU5OuzcRo0ntPiKZxoh6
CD6fZ0bfWfCmL6157ONENPqPbkeZP3m+rx8MdRl8l1C/bvLe0PFx8pAtfYSaTeMqp2Dixs0uxUUn
85G80ZT/G81W4k1+YO+pv5DgXTjhXeJS/KpwNvXFxxbs+k+yoB8JWZ+8X4YniMbhz506msa6txfX
19ZkErTr14HopmLxy+skVhVV8I6HqD2aHXL1dICphPR1i29OdTtUj0NK/ID/vhB00M6mAOhOO5Zh
/XUpSavMGdVoxkzzBAkBA+9QA8Kw+L6OKVjoVtLi8tFvsAnBX6dlA8SCAODwTKWYGx3M81mCwzbr
khU67Ey+jelz/W2lZQgWD/i/FyW3krAK5HCNFMW9WpCOtvbPvmdXYKfM+UiaN8kO03eIH0s+waaf
3UDMiUTEmPWtO6ZH3PB9RRO3qAf6ne6CIk0tORkiAa/nYA3UyyyhLfrYLfMIda03eNFrJeNQ69tL
nnd80ydjQWbuCCsYtu7qQDuaLmRe3bSyC63TouP5UxUPRD/8TG/jaoYv2wT0RlLh1fLYt81RT0tL
MhBHJSWPir80ww4q5XEWARHhzJPM3aULZSLDwWP9Nd++8R1yAU5bhAisMpj3iKpwxKbeZaKju5OD
nb+qrY5luHZRW/pWyxrdoqtnU9dkcKS4is5r/JDMV760hu5dhQ5UPiHgjXjXse0V2F+sNTqC8SBk
uo4vGe3CgnR+mBYieI9L9eXdnQWaMSSZdtT2GdkiAw2CDKjLfSL/0YaDYykUwH12piIIhFmZZPQJ
iiRy14dd1KLZMBqVxwAZHCsZZDXYixg4djbCIHqXWxtA7nwIdko0A0b8tDGMIzbAi7v8+s15IUsM
oCS+Tv+sPG7yh9kePtEmiQ5SJ5L/w94DNBbk2spD/+rnXQ6FZEjC/Tp7XEuBE6qn/YboEMWw3otv
nNTWBVQTvph8XsgOPfk7pyt8NYEu9Rwjs+eItbt8HzbPm9gT2b8sll6/SZlr7ddKBg/aMmzpyvu9
Ut7QmyGRB2ltpBCiya7yTZHbmpvIduNxnQRGjh+tKrS0pTviOo4Z95eFOI/8xhg5BXMi+R/9PGPT
lwOWB6Eo6Xe/wSWUvLB6z2rrdxqdZSQLRK0MWdHwTk/bQ4jw0yT17LAUdVKJYiKAoBAIIAiUa4iG
4g6LJ85uZVD/JMIC53mSlTHvZYUVw9KM5C7YChjLTITqT4FbEXvw8W6ASJ0FBoR6/4IJcozd2Fv1
/eLlK/ooLPdYeub/Oel8qObOUhy19FkZOzbDUu1lCePDO+vok5v4uFXcLePB2pfanr+2qjS5vwx8
nDORhLJP+8C8evJOcL7pshZ1tQGvIX6ylMP1JAvJMSwbWT1uEH7taxC8rYUhFOwXfCpXYsOhbqf1
WV7hAwnupOvqNPZZBfxru1+Ablh+Pq1xP+GO71kYN8prTLwjjeF2w8O+bjsYC6VhqGaqr+2bxgqE
kQpqRXsDszOxTAoe5beTm1fBbMqhtDDIScDya9f2stuTmdtUsTADvNrH58D98SX8UNQFdEpuFBTJ
uwUM1SmmyDNDCc71/luilCPaDQu+3BP+EjXzH8BSxYxyso0dcfuCUnMnrcFmVj8UOM04f6v9ghIO
EvE13JZLtLtimGanmB/ZH181Vram7YF8fl6JQdEbaJyh5Gt6h5a6iD+TtQQQ0Yjmz8Z7KyalKw/1
UY7OdOPK4Iqs/H17ohm0AzbRi/O3Jhyy+627krZPRmG2pnDfR5C7NN13/hbyM4spyODyTjATyELo
XpdElStBHV60pvw1VCdHClwk/vW9B5N37DlxvjMJNXp9HkwoUb1RqF/l6SsP3QK1ppvdg1DoFy3e
V0XzgMOmrWO+EJwMsZktAJeIgHYci/IIvFOIpSc0wfAVS+FUjmJrj/VMlUiKbQ1DRSJu37YQRJb/
NVlWbFaYXdZKpXRbZNPK/HEz6oZDI+6CkMr9OZ+8Dv6amsj4mxsLyKHPZXdkeq3DhPTZzYZ9nt3h
x6/c+YpAlACr4FiZ13YC213UcJiq0UEzpwbvTtks3dqgRBuZxXMUo3MuWfHQrggQO80eHT8NbAl1
z1HqAzQuX/CzmhyQLWQQquQYJESsbGs+UjsAYK8d92TQrxl9yWdtTWvNNRUEh75tyw8jQsPxvkub
b4XdevrK6uEg3Xt1qBqt5Gs7PlW1EtbYD8lA9zx1/7qMtYdemgu8aubcc4SdxMr0BOhku2YjZSOX
YFEPj74BCBsGThuc0VKbjNIWmA2Ay7VShp9R5YL2Sw4jZ0WzVhTfbCQl7prTRxa85JOD4oTzi2h3
Na48nzWOsjmrLwoNFXbRX+F5pRsTPcimvCmNjOhswc4E7TiBhEjoSkhKqNvmK2+iFQY72N3AXmov
pIDG/z2odHeRxSIP1BJtzEx8yEVJcEhAH+tFoOvC8HFJP1Tl8j4Yf/dRcJLWt0tjRFUj/jZY56Uq
sRsEFOwfGUMfDKag0l3bkzMy4L8XRIECsBGeeiaOdQkJcwFc086xp1Z1NTC7cIGn5k2hPVX7eTu+
+CGDTCmvKgYT0tL6UxlRoF6jwP6cIf2Q+GsDx1Lp+P8f+LBuMkc0GKxFUMzEC9JrtmZjR/fSA0L/
eVsoJFlmAsG5lZKJ1a7q03tW0K3NiGBCk359mII12FC8UvekBwFx+0dcV6hDe+NwkkfLEeudk3Tc
ITROto8qkSuLCxNeXsth8wWQnCrc17drNJb1Mle6XFM7ABeHopyILGnH4Ve6mQDmghlkolDAmoqk
PGINNEy2XNMPyIzqr2QGjWyk2M1ilWMF5pd0fQDufEuKFXuFjfXQFHrNNCi8nXk9gDtAJW/9hqFe
m6bK34MjDlqCT528pibr5XTOBQClQwyMlFErOL4eN+btD++ExRsRPN40Y5A6/xNkjCgENHErl8pN
MTfLMEk9x8tP8TwY8DSzTy/u6LjxuwlevLgW3wHsdVcNumsvLTjNs3pXMzC+cPvpqmCC55LEjVcq
YhRPmVapPLgkusPU1PL7islevEEH8bJM7TnkYxkKz5mOGdLLlPtGiAiT1YivK6fFytCDi81OK4qz
0zAMcZ8fhDhLbBECPgfZ0auSVMumz8rACMP8Uj45gHcJGDYZs+x/Wz2mhCgkfYViY+dBcLURuFyJ
AcK5ylFglPKsnr5IptUz44pEw2LuRmij2Bn9IrukiyoVhyXYsue+TO+6HQWC3VQm9ZP6N+r/rylC
aOwkJOBYItnqMVYSxgaXp/26QTwxXmme33yTKE5pZUv9Eb6Zeb2mzboBRQ6oHLpvNio1WgcP2kmh
PdDB+lmPorgJqzAApL291UMkyK/bw1gQErFzfYtOFAVmO6U2ObjurHn/FHaD0hFqv9LfX+W44Yun
umdMwemCXrqdgJocR8irvIK3LeRme6QZGfQvsihxw9Qc5ok7KsoRxtuFG/DzIupjXiJLcyEp+6Bk
K8f84pwLre1tnXuQ4TEyPTWO+tJXyZDeQiWjAANtmNcNhxq2h/v3yEfOX6DsQNxvyFnf9fQrkr6u
DfaEAWxQW0cMnb6RrA2JQru9+Rl0wr+JNVJDSTXxPzkQ3OIvvS1a8aTwWT/fQUyhCwr+P2egs4yQ
/F35uBz4fWtM3MSX3KPqr1Csle3Csm2CEPVUvTE2l+eMs3P43ve7zI2YXAFxvN8oaaQHM0xTp95Y
xkL1u18vYU22MMYhvs23w19pVJFbmRma7hm5Qkg8WGSojxKi+JeOGBLml8CMD1i7eykYVVXnZuz8
Doj6p5lhM9609wuzoeshoqzdYpBSTuoXogGqh+56nv8W8BNgBkWvcbm2bT/5vGACvKEf3HbU2XMZ
P746rnhz3eLU1guhCavl3bYQB8pUO8MQMuWHzfstO5HmapznlPEWEUkoidO5eiNCwjYkH4AZ61uX
NmMs6Xd9BX5HyQ6ubvNHfGJNBrIv4p1pQg2OQQzzEWN0Swd0mcFgDLr9DmVNVZNld+imIyW6RoPc
XIuRzxmLFy1Yam4hXGJu579yME2mHtjQzsUq1kjp3QBDd4uU02u3FJe0JkhZzC80zVFh8BBznOXd
cRdup8lI141oOaYmdsYrlLg+9W6J0aFlEdtOgWxAIkd5aWH1AM22Splq7MdKx52YuUfdy+PXncj5
HxccSYYVASAo8UCF1BXLECbgtTB5eKn+t8Wi2TnFmIxnZSdSh0eyppWOR168RihdCbZbiCz7bNo7
0Lt5gJNRof1+2qqSqev+TLOCQG3AxCGn5BKHP1QI9CwcRYbYl6qqrhcQIzPTVFNDbkb2oPjDR3Xv
wWaTb2qoiD421T3gxSU5yXHvjpPHcKidHT6IgGqB5b/hTW1Vvk8Y6RWNZ7a0WxFf83du9e09edO4
LOQ0Q5Qp6ZKcdhQgYLlWnvNHuo87aBMzSGUGlsfFweAArrwT8YS+YkHnKa11a1q1+VAFAW4w/jJg
Dko+0AC0SO6uLxl8FSqDkTs073dlTkFxOl3HBTzJk1k2vzzOaGq9U7VTI6e+vuvzB5/KIRPdtpi5
whWvE/rXehyuMcvT3BlWmIPNvCVUIsTCCOKwmmL5fQUFwpk/Jxv+YQ4JGQQJkOVoyZUiY2DXMyX6
oxsocwgmwoD/epPRlxHvKFyqSK+q4FLdwLMprQwVgf9E1bHqS0EJQQPpzr+mxOrLTUBnP4kwKv5d
G5Gsz6bQlFviIuy25hLuQRe259a1cxY1oe4mIcqNPOwvCYRatax2j4p/vtjwL8Gt1rZITpcyl/B6
fPbOPZFTz6K0IlXtYgVf/17nnubc1GpUd19lfHaSku+gjlIaQIkIAykBAduX7NLhZT6JJluGAYtC
L5+PGnzPVYrPpoeiyNrydOQRGddOf5CElZwg6v/YXLisudp8+AidWMiLJ1v4E1EJf+B3UrCibbHu
9H546zo8ZpWvho79rpk7gQaLx6/XP/oz/OdnyHZdBhfqe1LH5OoMJGZV6Q+sO5YbMzBL9ssTbUve
OPOGBboM5APkuDE2bOmLDBh3lgSnwe17hK0q3G7CuToHudBZZjTXTD6TEuv7cxjL7uf5OmxO8P6p
uzAZvKDyZRQ9+N0jkMDLQJbmfOi7m75CF7GukUX+DgRFrc+IrNFHI9BBPG3WIYLHwPV4ZF6AO7U4
E/FPQVSYZGUSIwWVNIMeKAIVVtfVgqEKErre7WtTq4u4ocfAVejMQ/sIlrSCDnzGkQ3vNiKGnSxm
K4NfJug+7xEdDYozyKxlmFPM6IDWtQMCkRBJCRn6O7raBIkVEdX293ye8ch2vJ7OGUo4SLRzDyZi
yVbDBPWtGYt9gUm38ZFzLEbv5N93zWkhS9L8kcERu5SD/igt4nounxyegGlMj6w44dO75VdPLPlg
6lP6lYpxrjNTtsIM5T3+b5p9M0So8/bO+XjAM6g9eEoC0e1Qb0Ugh95aCfN01OQgHvhVdGWBa1hU
+TsQwxa4SF+qmUaxXR8PSyggW+3a71wRqw+o+fDQiPybsSZaEWVv3VJw3wX4kk1voC/uk/mBMh+s
UJPo+GI00xhGxWlkHbacWZerLatORs0ykcRw6iln0viKCySv97yrbhDIi88N4WGtaV6I1HYWT2io
t6EJ9iATktawDvCQBpa4wsn8OPYEWulP2v9pZZvmNXM04uLpoKUP/CqCN1U1CXnAyY1Ws7928wcO
Vlw0/Aft1kWtBjOhABbxiCUgv/sU1tIUBceSk0dZTFYHbx60+78khoWHqYobR98vzcG18g9kQq3U
0iQGEW1okwx+4nDBISoT0XumreVaCu2tDql8/lE14rrJIUtvxw0sRPBlLYngqqjAwYePav7s8GeC
E4f+6C0k3BrJxx0Z7nPvF00ubqkEISLZvWFmuXpIBtRdyqu6RXMOBY1Py55KBM5hrQ0sySDSbjjq
kquUEV3u2ukUAyROBOgALzC7FTy/si0iq1r+2oX2L824MeKvv3jTSxNWu4QxMDZyagOz8wnIslr6
TwN95jP/87K2ePH/faZSp+e5mIdqgDSfNiRdkaaP4POCfL48rhvVo9b1ejN3XnwsRWQ70mIZAYhB
K3XNpTK6jC+KAFwGIMq0BExbwPANCWhldy2CZhWW8VE/0gYAZCeDoGW2RPQeiOE4kndvLePN8o4q
YsbNl/1lsR/nibVEBCEAVElxnMk/WgHk1suiGaIipSBXq/5I/F4ZsXu/QYAEKc1i7W+khhF50mB5
PlsskSm5Qt05HZinU8kr5Ogj1sWQ1H/2zBN5k0ZgrQ01BnIuZjOY6zHJsrsTk+D+nf1D8zFsSjPH
XyMQq1eJgHACj3Qj8TdViUZ/VTDGgE+WCujzmWCnd0euDwMQ0ydCkl2Y3x6RRV7zJ5ato2JQj74d
E+SUwD78xPYV3DLgBGxIKxoxW1y0WUT/oE9E7lSI21F8IgGcNPpe9Hh12xxhYneewzTfAmNaj99U
cf7vRIQW1z2KtAtbTYVqD68VX9fkfKDgo7F4M3sg0vOKnpFOl7YsMyaI8O/AVHp6ZCo4Qao3pjWs
qqJizN+KL0dlqQAYXYN1uhv0zxCscLk35pl27Sg/+Jo8ByL/3J5dcb0oC83RHX+58xoZz5Z3ynww
SaP7px3uijB/JXyf8TUKNqPvGOBkcOm1r176B2V0KnbRiSYoRCij5dinZLc6fXJUS8adsVtJ3WDf
QKp24S+URHqIiZmEzVQUJ3ikN14ps+9gmfr1W87lljog/J+yTr0a7eLgYFqrHen/7qm92lwMR4Gn
f7nKbwG70d2ISTtFmAyTa1a0fvWg4Csf3PD7rrMKo42V++wboWkKDnEqoulYftqbNOZP08+ZPrGJ
RWwRtkVNiK/PKXz74facIb6GJFnksNuzN9O7y3+qg77spiaNkfiQ15YizF38Y8Jmk/P1HpIG32eE
WTLgCPJ4a+7bmz55DSa8KClBf7fvmWoCcTjWrYMrnzN7hIgk76Rw/DQTenkC0RvMobezX9Ogm0we
IKgxELVcsfHXBX3d5AuBheS3pFtrbClftFW8rnnEquhPKvPDTtBgXsQrpHFx7Kvia86y6rALs2NM
Meb6wK3T3WVTO+mkG53cK/VTqf391Ajv9xMfXgWbTeBLA5Wq1rxlKPdAjVU5GqiND1Uz3GCVyl1Z
9/UDA/YBIhQxGzWKbGcaZP3D+Q2XRBE779ySXbv2JcdQwnNB0Ubbz9erS36lbmzCjnbrMQIF+9Mc
ZFN5chtKy70KaUPenhH7sukTTaVWPVJIoN6bjp02IbM37BcwjzheWEpgzPES2dy1247yh2yQCcGc
lMXE408xncXW9EOGgW25/Ph/l+e4WLgtaNAlkHfZ75NqrHbITXXXcrZZI8mr3AKnonl5FdNFmp1a
bkR7duAthsChViBLI+8NBXo4aSp9B3tsczPwr6xZCL88PIVJv2crLyjisSod7dHC7Q6hX+N2h9ot
9bMI0BGDVWsuibJPy8uD31n4BTW9+bE9+n/vVmZXIXenKOIWyZfBipXVSAlDXb98E6a/uKI2kZRV
JpWiRfBSZ6iMpii/gAE6b6VqOwfhYtxvojB/tGy8Cn8R2UGdFEsD56VKQ269fPB3tiLc1UGHyqAp
3iDZD7Mcc2hmNV1P4/NQLHx/RO6x62cMw5e1JjFfs+ZNpzfUS5BlRyoY1ytGQNl3SlGz1+pvY1/1
rG0ENMYXjqYNKOFhBElk/8Ms79hNgjbtzzfVHyXw6RL+eE6RVkV/EZB9wxtG+CSOsk1QOYjzV1nB
LV+6GLf0cKFufeSuIwwplPHj0oFpdJqvyTNulCUCjXR1OVTw1EotBVjpTSv15VHSblBhxgYfx7wP
vEE4mj7j7rUs62bJxa8Nbemdb1MQDCD/NKPo8okLsAoQPbUHHmHIn5NW44RK994uIqckx0OPTJRe
ikdRlR9aAPEuxTAw4kZ85Jx+k7WP57XKbFpR67T13Qe9ZnwnxKh2iVmqsJIxKY2TFRbNFAqvFbAI
y+pQwUy3mafz0B4KIUkGvDCKSvMwxRBZDU/bkTxQP7Ti6Tts2Jh8b+CGoopiqsTWfzVUeVw1rMl/
9daD7YPflsmPFQaCsh+EP0imw41BGbHXR4Ym3pxIinhyFVpzHiW3KkX4VxDMu92NoLJ+6qCSTDkB
TxqyV6r5HLmWHCmPA7lGUP3XGIAZTLCD6ikfErpT84v0jJgRe4NeX2X809u3os5vcpubLHIGIBba
5Z+d0+Nr6KbsLB8gelfqqtWquOUvevr67MKwzCT0lwiDfVnsytatd20u2X7zeWKV9RKcnAMSrfwz
yTcAEOMTnW+DBmFeCPR/nuGPWt63PlC6p2uGx7HLPUaPX4Tm0zQgqD9GgNUX8RPzVUaML7PwCUVq
uz69OeCw+ofVm8Spt59AwJDS7ff07l7yXpS3gtVNgt14IWUYoAwJ0qPQ3mJYmVqtDbv9i7/EAwVb
CmxvTw5D39oyzLUwJqm7SMsUGMCHjdLJsaG6UvchVgC8KJxLbziq/wwfGgkyFEy6l9dhs7ER7uNn
5yTuEF0aEtgeNEhFWxHcOOLcL2U+sTmbBHHPyhtM0C47Nc6Vy8jJtsHylSagPg0+FelnETohyq/t
WLdwdup52Y0bo6mbhJMhmpy+C/hz8mU0q0PG0FeO8mGH/h7UYGnMEj/cF4i3J9Tgf56H+FwctoRA
xzM4ukC8lKcl9YRoTgUsurUHmFEenn/Pe7xxtL2pmFBJuqdXLvtk9PnAESXiv0DucM6DJJ/oC9t2
8y2g3Ek9zDJeDnoqif/F8AyimtcxAZ5SO61bJtlB9bKa+SHJb1/QVhYZ5agXzJAzlLycuZstaQNR
3U3WRkaGYJc0rcgKrg+V5+XatfLg/+8fB3z1Jbt5OFqVSn5OMt1qpjgGHB180GZ/xcEGYMhrqvEC
YSELD2yrqBJ2ZH6f4y4kFQepFxuHymDpPH6E2ds9T7ebtz9WGXFmmMt6uYzRPinF7BByhO8sRh+9
P4v3GRZnNXLmjP4HJMJfXONn2Phczh0l14DQ5wBEmMUs6SLr6UdNcoVcsJrcX5X4O2J7D8iVTVfL
hS8BVrrxXwU7zXQkx/adE5hN3HV8mglESm85/jC3OLqGm9jV6CEU3lPyuHQxPZH6UC4ywlTrqsLA
j3qCGx4ycYqMmwzVYYFoITdLq8b+HUTBwuz7m/UxV4i7BLhTLwBIjRkmBcVD5NwPyVZT2mlRlngM
cKyPQriDrnDC+Bsl25nu0lrfsr+EF4VEjczLSkGk8W+NA6aABL4M3Ss64721rrEth2D9lyHrJjl/
wCB1XZsS6ByGlp7O/6mrZqG1ee1kYiPvU3ZI/74qRIPkFHzExWfqL4inea7fK8kJeRSwhm7ZLgLi
x8A4Zvgnz+q50KQ6hToZKwJQZByjenBbmQuqwnpSMlVgNmG2Ee7b9TM6ARIics9LFIIKj7gsWYTU
0C/7fvr7XcKRSjpdzJxLlT6QLYGD/CN5Gzgp7U+FL919cNEfR2bMDulOoTHLqv5d50Qa4KRW3IcE
eSBeySgdBpPuqBmpJrPeSkkUs2LhGKCYwluWJj02Ov/xPkx2uQLH1RXKlrRnajK8Otwp37/TAvkV
NSZ9jaQ4l/nCTOBqNX3VsEC8EpEOqc4pnxzO24VRubzOgktqy6acq/qxgtvxhW6YDDnKTfuRBixM
956+cS5g5cchB+m05YCTaDKB0rSWzjLTtwVv1GJ0I9O2kwRcSX0Hv+RnefU/IMZSR4VIo1KWFytH
gyAVdU1GjTIKjynGF/tnMlVQMz3zSrci+YQUFntZWqAWTJ8BisTy4Nzs+rtYRgnd3sVTljNwkCPx
CtiHj1ZWi0/LvLoJ9EdjfcsTEStAhTFV9C/CsBZAS29j8oqZewFJSBdFnZdlXhSPELekKfwMcVxn
9jGRh+Z5SHlwE69I6GPAO9rFINI0ghVcDvyPmUPSFUEbBqf044JrqC4M9JtEdzRpJtZwt+3mJpQv
A6waJvnNPvH8lSKeBUwPC511EMC5JhKH4KoBv/9nua39lXqvfSzOZ7doLSejfqN72boocZ3ypcn0
eb4seCdXRoW+mvi+VTL6L7LF3Lm15+0ufWh/h5xuV5v7l1wDMSJW4X5IIoA0dzJdv3/Zuoi6BI7U
RP1tTXyInhOtZxbQALgW+Zk1PXoPrgLpYMyN9Gk7vxTYlrtQlcIZvGfaO8fDT62ouSgVDFUN8ykF
BpbUDZiLQSm0c5b+SNZ2iY30ZgHUyYAL1pYzZG6R6CqJ3CCdR4ZefSzjykK0yJaj8/uWsWjwSs5+
u/xeMmdiKELYUn69viwVzc7e03JHdLmiU4+XHYaaT7wJTKH5SbyUHqrlAV4qKWmg1Rsidj4U890h
GLi8cdL55TD7i+4HEiIp9K5XS+TZRPVWuNCRh7hX4dwRP/esCglPWowUmUW1gjKI9xOF0uMUkB4c
JwF1AnttJqrnvqtKKvkuQ1FY77MQhUicbJFPxfKWgXDpbsJURTajrwIN9UIzvVn22qhqHKc8ulrT
4GaHTz2eb6ZhL1mRck16XiACVLcA+oc0eoUBwCGffcBQ/4uo5tr/tgku3cVaduZhQkBNUm8TMmZ4
+FCgS3XkE0WOgydATeBqh/HeHLKJZchzqr+4G1eR8Kn3kreAAdrv9QP2AdALpkxQoP8zFZO6p+W3
6gJHhe1qTweroRL7MjfPAucyZK1XauUk9D0JfzWNJ1lN/3EVpAjzLL+Nv09Pelnd0GeU33PzKbRe
2qlptHYcpC0dcGhaFQe2brmAOGgGQOGdDDHl4ntIDUR6yeJUIomwkjV9Q2Yvv+bNRBPa7ikEPpUt
+cdODuqPL082Hs9/aNg4oCN9QnKywH0/ocPwOdWA74u4Oo75ifoQ7rf2HD8r2hF/9v45O0ENW3H4
V7ommnO4ur2PbmW/lQHIyRO0kqiNbfupwUjh0rIUvFEc8FzplRs8BpciVbkyjdWdIFHIEZZZmIOP
b+Z6UreIfTgQNcL6vvyMdO1NN8NP3wz2QW2igeggMVWGDMtgaiOKYbZqNUA/qF/fQNYSBDYVazIK
2sGy3mSaIEEa8qDoXBr4RKDuRuDqwB3qGzam752FfzFMWRl5CW6dXMC9AVod+b0Eqi9z4sHQNg2A
XtaWT+cNuCEkQx+dTH6e81bBluG4LwqjvErkRGTBR9xOgmhgOmgfCTQVzOmOtIR342JYXPF2WGD8
XKh7qHdWAZes6dWgscPEkF/GiI4UVRi/06dflMSmDgOkv8pnFjDnSRSDWnLmggZ3cpIPqdIhJthw
0mooc8Tr38mEUHbsCxhIP7hUiiN7m0eDZraV3JRVpSkj5YIfk55oYUyA+SxcXKJk/Km2Sl/AxVIU
oBtUjgicYa/hv+ZNBB0Ie6qkCaqa0ecnflpy11nIkXEDYbrbQ/dZnWzxuc9Ec33Ynynnk9cH1KHH
aF0DvD342YF5o6aJ2oibmOzKaxvPdd9P7UK9AH2Ep4VSsLT1NG2e3AjosXbhrWuj5E72cHTc/uV4
ay9qu4xW2vzaWvZ0rR6Sr+5Al4cPmhll9/TzU9bPC83TXBgqOKFroG6E5D23P9anbgJ1j3IZ2Tn5
dQYjr5NajQGAkWtDvc1En4GQOosMQweJAQ6BKOqn+diS8oODnazY1NbsaQfpVYwI4IzaLYWMctMk
C7WMeqLyhmxouiJlRfpXbN3XXNm1KZ4T9Gj5xvIDUP0hDAXvqFnwJt/CI+oASJCvhSVHKyWFX/KS
gbYUbVbMxDKbAy71EPWCKkgA/fk+3yf83PaYeJn7KMteXjHXr2tbCOWSlgR5HQkEAuRFjz3dK6Vu
GSz5nzuxZlAIOJ9UJ3n+ZcRHbqB34LNnqFpvC9iOX9BEu1hAoe/Et+Az6JtZ0r1zOUNg4/+k+g3B
6749zZWZ0R8rBYNKBOyYISg3q2yycd/xjDroFwS9Gv8hBB9sgE344galC4ZIZjRzCqZFNBA+SCzH
jwWkSq+IiBoPi8qPdwa6K8uhHWq2emsO8wdaUs40BUfEulWkCRGbDQVqfYihHycxjq5PCZ2pk/Nt
Z8IaZ7K+Ume5KXqtyCmuI3D8TGeEL99RpluCNW/xw6swkRj4vm/gIHb2kRZGFRgeNDdAUukXXnGi
Hl5QLEweWsSzHYgFQvlLHZJ+FlXtY/bd8mcqzykSTIP3y5L0dok/uAIM3qRqEoOR22YXVVFfTAHd
k/tdFcgkP6Jrvi0s6ImVo8rh3aKuACQh6XvxvixM8mAj3EAfdUy7a9G5KPG0/R7yQ437L2vxs4cr
AdLC642CPsPzy/xNJoHgCoj+kSEVxnyYtNINTMoL+Lu1CTuNhLotdQRBLZAjaz5Xouj5/N1MiD+0
FIR6TrUz2vnKr069oCb+hy4lWpDt+686vpkk+O26g+bUgkJsFedgYJE1lMpx7ANk8t3V0tyXKL8+
memFrpjJMoiQGmSscv2NAWmvlKtAaUMmMVYuYTisS1OJc23kKnRW/cyDyazskfzrlryFFXZ+z0uN
O8Ld030AIDmZu4SgfmWrvgldCPDChA6wA5oQ466wOdYb1V2OIrgRHU7iySJ2k0ZJkYOEV0u+aPmI
6KBTW7TuiJATO2kwArTZ2KesCpeV5ZY0meGI/zvEDCpErOdG/Au/YfY+Lhjwlv6si+UnUYAFaEEW
+2Hwcsrh6rIZ54msY/Jjcr2y8m4Up5cc5tyfDZek0vOyQ8Nkij+XDFCTZ1rq15wQOm1bDNbpEUNw
uQ6ZBTpwKrEZayLwlQca/wJMkBKG0mpSEPvgak/cD3aJQ6iPwyPXwdkI943vHWJBfQRTPA4XaddT
xWtpMVAtA3qk8qI8/pIqrpafu3br+Ea4QCtVWmNnch5WgU48PvlhvhR/BMOURhECXTjBIq+aKzjp
XRnrtUYR+dcrg8b2kSIsVRQKPlYruR+GGRSdbbGGozt3jQoGILZYv8SKWjA6H170foyfGgOvcVba
+RMD0UtJ2s9pk+pbMe65h8YqmI0D1F/In2U6axPUVxBgC1g7B1QuUeCQeFUswMeSI6yTA1xzbgZO
yyixeb3Oj0GQmguxwL5PBKy3bM2TyPkknsHQ/2Eyo9ZsGD1PdwIvf/oKpvSXBoAoIJ5iwuzmxy/z
HfHD4tkLolF2RW4gG4uTR9t/hO/PTcffbezAV0dlH81gYV6OXVhxfW2TKI6QaOBPEAagZVrhCvr2
wxshtg3sVzdCZFS/pZq/IdsMwS+mBWV48k9+Mg8GRwv0edfRd4Hs53x39xd+yiy/0yVNFIfvhYFB
5TO4n+7jj48oyhkSMiHDIab5CjwqoT4gpf/FnVnox6OGoOKVaTr/+ThScc7+L0fQXdMneXeWfwTj
7/QRBaCzyEUnlPyOwrtrJZZAbX3EqvKjMaQ4dfdf12b0iuf0THTviggUEvvKM9OjfonzIa3ldTjo
dqJoEvHl+iCpAOu5KzZPWJpO3FMM12PNbNObbuUJGHSyY1MV10osodTeQyUJl9KVYY+dzMeJQSxN
KAZp4hNCsxaZhoYpfqT6zuA+m2zUE5BFvnLmrPEx8shD9bARQmuy6OG2U4S7WCmZKouKder+aT0S
q9HJh7G5jzRtWcdK8+XJMBvlAHcTMJaRCJu7QtI9STS/gHUFUlG/DjxU5Fj2U72YHSRkU5zhig9v
8jR8nXsyNx4RqthCnPcQ2IkRB9X153vZNxIgxoXdgQc7k3FBuZ7Tx75pAC7J+7FvidBhROmhMM0b
HflicAzjjsl7dq8DlVL9j9A44dKOyxb35pu2AL/XkIBGYOpDZIffhksEPHvcx7oYot3KdwYP/0Cz
V0fsdigqp6VKdH7WrMZltnlbYyGZJQI/cOQgfXYK60UB/8fyT+T7YdxdPnitSmhLDKxBfifEu4tU
IyncuKEc7k+YIeonQk9IV7x8aan6fv3OozDZgWJrZwajlOeSI4bQdjxpJveaxsuFd6BOwsybD8IZ
NPGWPEhBBulDKW8QeQ5l+A58etTgltngS9lH3i1o8z1hT1XHI5zHLox1+hDWgvQCvTvskyGrNM4u
wdOkTX0Zg0mJ5cjwflxK9UTQW6pZVZq6n5nUgeEInyQiK2WCQy288/HV+kiDneMnhDqDFVmJkjB3
oGZwsyjIyN0u4uyY8XBL6J1OaGqRVG+jjQlRpP+Eoh3tR+DN1m1ZAj2NN/u9HKOE+OcAwYpYYjNr
usBSNgFJYGFTMaUhUXZL3Sboq1G9RZLFg4NcAKC9fjFmuh9Kc4VN5MVWsDAcV2Xwvf5s+1UPBZtJ
3uYLglqcSljM+Hbn7cq7nvokQ4uTt/1zXNCaWPR+8VuqCuVdRY5NrJAX36SHy7rBJa8eKOJaXEAu
EBHhrETgiRNKlXifH1SyaQfFsHQ0bsvWkHNodNRvledR1rXaxK4fzJbzXuS+oFmjtPc0w7WJfGgr
m+r+ZZ3WU6TEUWv7mA6FbZqYK3SqYNkwXNMbE1SrTvAhvJmg189VJbTs4lExNKhbCQuXGQ6aBt0v
wwNLswI4xqet1Xuuvf/+g6fd8pOPNeWK5OFgS0ovnL2UTdI1DEz7Qo3Rf/S/dvHxNimCVCIBUEhu
Vsr0bjwYTXz7MAO6n+2pUXfn7nXu+zrXgVX5zpI/r2sUROqAkiU5TB4+SkCp7HF7QgMEadZXsAQ2
acqzzCd7O1XarfcHj4dyqLg9SwXjIB5jvMNO9Hqbh3gf/mfzrm7Gr40T+f01xiiyq2tH0DVhGIuY
eFOe6YXwyuOftUdgGvPzZ8aopWbmSuKSW1gE8K+KHNxdQu69ViVqOXlNtGF1E6XOGknEnRCUL6E1
f5ttsWPxr2W5I43g6S+Kscin30toFLOvGs6ygM+wMWsRzYhDOjKas2nX+JyZZo5cdfDUwIasqYd5
qlUNxYvJoN36NX8MvhyRQOxc4P37epUgHWieiRVtwWjGG0sVT4c8KHWAvqJ5LwaXgS/EDvOQnDWo
SYvWTqw0l/16qWiG3aVA/sCfNPrPeuCuEQ0BPaZlGZ9USMxy+E84NBSms5wEub8IFXQk83Nc9n6H
0YgiGOd6hx9PtZBppf73aIiSRlGyS7HfEtOFcHayMJBWgZSX7oPdTuP/p9lvWZ6pUIAbbTKesaDF
0uq/mWrbQGV2lMkwJQGOs3Pnx8MgM/0VwzHMIQhceXK/qpDjZI/j1v2UyI1Q5931/fPbnZjgG6zF
EY59JtiDpw6vbY5LsOc6OE1RuyWSi1qfp4yd2qcsu7HlmzvkpMWL3qajrejHIGxyPmFBwWGHQH3e
Q4BMmLHoYqHWuZwlOvxtfTWxtjhvVUKurPpIadZxHX/ZNY3nUNIxmE1GPDUnvbcULE3S+3Zzjxkh
MHmfN1YI5ggNIoJVQA1TOSTq28nvvFY9vH2DiSxJYgk9UjzVKEAXujrvjcgWzMAZZBhVtxj8vU7T
n8XSycUkKR4nmpYHt0EgKiqpsm1lQcrb8SlQ+YW7DRSpmPyHRgg0/I4Le0ZSV0F1FwwHAcwxUeDr
sQwQyYivFAemzPoSflk/mPqr6jOznZIwZC53Dogi/BxcE1fTvijvtFEpq+vrLXov4K6F6lQYuG5X
dg1Qq2e5HxkNwX9hg8EAGUJ8tpr1gDv8/RP4NguLxPQA4Eab1MXzh7kpnLXPSCDCr8HkV1vMMAqG
XBXSz/u2EhA+U3O/i/re1CNqkaYNdQ26+E9XWE9tz+BWmGEGLwWa/svWSvr8yINBM3xxqMrp30Nd
t7mHmb9ryiY9G43SL4rulYXnjzcw1JPVPNjUZqpOZyooDxRe5BKF87LxC4SnyodlfpD8ZKHuD3Uv
Lobr2i+8YjPClc17yPMYO2ANto238ydmqtil8msVXzXS4uBH1iJVTRx9UEV2lM1s9jeiWIXu/H/Y
DesEmDpUUfg9Emc8rBLuisNoLF8iSdY2fuIpdKNdVMQSbw05+TLhhOLuVrYI52XTQCi6BuyqlVYG
2jopynajaEtQ7E3IvKGK8t7gYfj49eDZeicupy+A/nWhsDY6da1GJF1sXhr4LDoLmnFntu9ejlDk
FAMAB5naVGxKbMbfbCb5UkSsVi9o2N1zQKB6oX0OabRu90DhNvSDI2jPjapNCmSEQW/l05Q7IL+j
MIPGIeSVr17NHhOsUYo1etVESaSs1UFNveAvOGmf7p4N6qqgmJe9sTjLE6XvaLlnRHmVNdIfbcG8
RfA4XVUg6AhMPgiRwJrnftMT/mo/DagoyWRg2pn+ey3Q/CdGLVbTn2X/I0vmNpqEcFDfuGAa276N
+M47wWz9jq1bdlo+QScrcd4f3zAFSdfdiuBKtzgMPt4XzmSrZ3yvZtEm1VOOLRda5P8UV5BDxT0q
prSqQKZz0LbJcP65ffDOi+YZf//nkCotiKZJHlVXzZA1VTLQhgjVJXEcP6/LxROq5HcqCYD4yq3W
nEE6hZU/hjHLLZ9G8zTDWtVhkP4j4MOSUkEmKVp1W4/9npbDSOj6qpfBQ6q/wkZN/vWtcw4XjuYR
38nEunmWqlGRvzAk7H33zrFTgFcBkUFNIdajO47tiOEHlLITdT2LUIE0fn75UbkDvgYOsO6iHZE5
FX/NfE0AX/CfzCTtz24qMI6YqbuWqezjN+/f0Enzu6JULGkrFuhTnm1VGqAmNR0k3I5Mrqzv44hX
LAKIL0nAB1YWP/fWVKz+93d2J96fBS1rbhP3r83DLAtZAS5Ihrd5DbGzliD1GjyjzxVXFbYumlm+
hQ7BOh7BihEU0mCuy0K+jdy2qS9CbPuK+Tf7cCquE/SpCkDsqK034vFMZiGsvAQEP835IXpdHmTZ
qdlrczhqR5w89Jc2AqJ08+Mvtie1IWXA6WFwcCyuJxfAi2Ujamv1wpzr7SVwQekkQzTqAyo92jCd
2Yw8ImMeropmlc13jyy/+Meb6sdcvn/Khy3g0tPDPWMZ19EYZU525VmZ0KqB/OfBZOw+oK/HtzpF
dbONbb5MEiQ1YLGgjeecbrTeQ1KFlZ2HWQ9o3JadVj9Az+Iu1vmkb63XUGUPqF01gmNJQ7AifNqr
1dhP6G/3G+2A9FHTI1Sc5IoAzWqHwM7h6eGFelW7goR56SGu7GCyGYlseVQWqHSxSUK1RM7blMg6
ZsxTwjDSQ/vZtFEt1iU32lq+w09iv93DYnLolBPhjUSkvCAfP5GDVil8jggF++N33cAS2ZfyBKmo
HnA85Aut1sIpyE27FuvRrjX7Ws/QG8D1U8DkcgiIIWcOu71yp+Kn1LiOxalTG2aO7g4tTP5kUpOu
d+S3Hi5lzW4pCiSjDNf9Wa26HbPpA8jbzyIRzupgocZzNSH4TUlCr0aC773eZ1cUDESUUOeyt14I
/txKUBahLo5MsvWnS2nsZ9kVMW7u9Z3TMLH+I44I8LhLEf37JX8Njelf1x1IoXH1JbS+KpUDHjDJ
//S92i7poRgdZn0dFkbF9wV0tzkA1TMboAbHf1bFe8DdA55oOdmQ15iAqh9ixGewXm/ieKQkYafL
yOCkimZTbhZ/KxcGHBcw2MhYrNsBV+SSjhDnIPlvE+43awRwNVfCbxAonN94D8JDL7w4sD/h5mOj
z48fxARYWNJqFjOLoZq2SjLmRwXLisRf/yc5OGxMDO091WLB0NvX4bw/WzypVBz+aLGMPYJpAbKr
HTwQAvQ8WsCu4j18D/d3jlNP2GnlWJqGRVLwRx/C+1+z1ks1t46SiHNBYCwPEk3DtwNTvBlTFsGy
XyCws3DD6H1o37JtNq3VCJjs4/6sg8K+6FlxeOLtUen54Sc3SlWu+IYFhTQ9mSAjp0NSVBKZQ03Z
+24x2Ow+uk08tdLcYKmTmfZC75vMlcfHnahUu2VBHs5synhYRZ9xXr+i0499YyNgeAuq+jdfQ3VP
BayIT7C67Ff7H9hnfJw72arDusYQ0IJNaSE68V9m67SAzJC5gRA96DNvTTUAvNt8pNAQ2O107oMq
8gxKqA4hI8IwtGtb2FTU7madfZG8fqzCSnr8qaEnn2cC5yrNz6WlK43jpWAkYPbn/2pFkWYMRgnm
makrVumiZQQM1rPKPvGVPDl8EAZWJhgUdYxSRo0QKbBksFCEdQYIO2LM+9uNHnTYNzMiQkCnzRdy
KfLHqHdcSmD+8R8BXJpWAJSokS/m5b+chOcVWwLJJtO1cIZ/3K3OFFNI/h7RogI5Plm46YzggQSm
L2jJyX4gfUUQlRUV3Hovig0frWUOdPMf3cdBXq++pTTZ0rhAvL3R5g5vcM2fJQr3H/vSrmPhy8it
eSLpivOop2oV7uoTNlN/DbS85lHGPlTAo2S0Sm4kANBbXMUzJx+cX/+Pg06MuxCsJ6ugRRAwQxRj
h1VkACI9TxAuckGNtIzXpuj6Nf4megm/UyPaNV7HPQyseAOrzz0LEb0640lyULPo4jiq/7nIk3OG
birT6GgbBGJ7FQicn5AloaTDYiHcTDJMZLE+kqM06jyxMR/qd9Tl66M++N/dg9ApexHAJNX7kZrB
MWhSH6djfHYGyPvhFQ==
`protect end_protected

